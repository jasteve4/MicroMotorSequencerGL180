VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO driver_core
  CLASS BLOCK ;
  FOREIGN driver_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 720.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 687.400 -4.800 688.520 2.400 ;
    END
  END clock
  PIN clock_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 706.440 -4.800 707.560 2.400 ;
    END
  END clock_a
  PIN col_select_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 573.160 -4.800 574.280 2.400 ;
    END
  END col_select_a[0]
  PIN col_select_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 592.200 -4.800 593.320 2.400 ;
    END
  END col_select_a[1]
  PIN col_select_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 611.240 -4.800 612.360 2.400 ;
    END
  END col_select_a[2]
  PIN col_select_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 630.280 -4.800 631.400 2.400 ;
    END
  END col_select_a[3]
  PIN col_select_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 649.320 -4.800 650.440 2.400 ;
    END
  END col_select_a[4]
  PIN col_select_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 668.360 -4.800 669.480 2.400 ;
    END
  END col_select_a[5]
  PIN data_in_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 59.080 -4.800 60.200 2.400 ;
    END
  END data_in_a[0]
  PIN data_in_a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 249.480 -4.800 250.600 2.400 ;
    END
  END data_in_a[10]
  PIN data_in_a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.520 -4.800 269.640 2.400 ;
    END
  END data_in_a[11]
  PIN data_in_a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 287.560 -4.800 288.680 2.400 ;
    END
  END data_in_a[12]
  PIN data_in_a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 306.600 -4.800 307.720 2.400 ;
    END
  END data_in_a[13]
  PIN data_in_a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 325.640 -4.800 326.760 2.400 ;
    END
  END data_in_a[14]
  PIN data_in_a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 344.680 -4.800 345.800 2.400 ;
    END
  END data_in_a[15]
  PIN data_in_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.120 -4.800 79.240 2.400 ;
    END
  END data_in_a[1]
  PIN data_in_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.160 -4.800 98.280 2.400 ;
    END
  END data_in_a[2]
  PIN data_in_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 116.200 -4.800 117.320 2.400 ;
    END
  END data_in_a[3]
  PIN data_in_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 135.240 -4.800 136.360 2.400 ;
    END
  END data_in_a[4]
  PIN data_in_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.280 -4.800 155.400 2.400 ;
    END
  END data_in_a[5]
  PIN data_in_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 173.320 -4.800 174.440 2.400 ;
    END
  END data_in_a[6]
  PIN data_in_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 192.360 -4.800 193.480 2.400 ;
    END
  END data_in_a[7]
  PIN data_in_a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.400 -4.800 212.520 2.400 ;
    END
  END data_in_a[8]
  PIN data_in_a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 230.440 -4.800 231.560 2.400 ;
    END
  END data_in_a[9]
  PIN driver_io[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 21.000 -4.800 22.120 2.400 ;
    END
  END driver_io[0]
  PIN driver_io[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.040 -4.800 41.160 2.400 ;
    END
  END driver_io[1]
  PIN inverter_select_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 877.800 -4.800 878.920 2.400 ;
    END
  END inverter_select_a
  PIN mem_address_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 363.720 -4.800 364.840 2.400 ;
    END
  END mem_address_a[0]
  PIN mem_address_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 382.760 -4.800 383.880 2.400 ;
    END
  END mem_address_a[1]
  PIN mem_address_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 401.800 -4.800 402.920 2.400 ;
    END
  END mem_address_a[2]
  PIN mem_address_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 420.840 -4.800 421.960 2.400 ;
    END
  END mem_address_a[3]
  PIN mem_address_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 439.880 -4.800 441.000 2.400 ;
    END
  END mem_address_a[4]
  PIN mem_address_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 458.920 -4.800 460.040 2.400 ;
    END
  END mem_address_a[5]
  PIN mem_address_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 477.960 -4.800 479.080 2.400 ;
    END
  END mem_address_a[6]
  PIN mem_address_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.000 -4.800 498.120 2.400 ;
    END
  END mem_address_a[7]
  PIN mem_address_a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 516.040 -4.800 517.160 2.400 ;
    END
  END mem_address_a[8]
  PIN mem_address_a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 535.080 -4.800 536.200 2.400 ;
    END
  END mem_address_a[9]
  PIN mem_write_n_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 554.120 -4.800 555.240 2.400 ;
    END
  END mem_write_n_a
  PIN output_active_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 858.760 -4.800 859.880 2.400 ;
    END
  END output_active_a
  PIN row_col_select_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 839.720 -4.800 840.840 2.400 ;
    END
  END row_col_select_a
  PIN row_select_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 725.480 -4.800 726.600 2.400 ;
    END
  END row_select_a[0]
  PIN row_select_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 744.520 -4.800 745.640 2.400 ;
    END
  END row_select_a[1]
  PIN row_select_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 763.560 -4.800 764.680 2.400 ;
    END
  END row_select_a[2]
  PIN row_select_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 782.600 -4.800 783.720 2.400 ;
    END
  END row_select_a[3]
  PIN row_select_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 801.640 -4.800 802.760 2.400 ;
    END
  END row_select_a[4]
  PIN row_select_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 820.680 -4.800 821.800 2.400 ;
    END
  END row_select_a[5]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 10.170 15.380 13.270 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 190.170 15.380 193.270 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 370.170 15.380 373.270 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 550.170 15.380 553.270 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 730.170 15.380 733.270 701.980 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 28.770 15.380 31.870 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 208.770 15.380 211.870 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 388.770 15.380 391.870 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 568.770 15.380 571.870 701.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 748.770 15.380 751.870 701.980 ;
    END
  END vssd1
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 893.200 701.980 ;
      LAYER Metal2 ;
        RECT 9.660 2.700 891.940 701.870 ;
        RECT 9.660 1.770 20.700 2.700 ;
        RECT 22.420 1.770 39.740 2.700 ;
        RECT 41.460 1.770 58.780 2.700 ;
        RECT 60.500 1.770 77.820 2.700 ;
        RECT 79.540 1.770 96.860 2.700 ;
        RECT 98.580 1.770 115.900 2.700 ;
        RECT 117.620 1.770 134.940 2.700 ;
        RECT 136.660 1.770 153.980 2.700 ;
        RECT 155.700 1.770 173.020 2.700 ;
        RECT 174.740 1.770 192.060 2.700 ;
        RECT 193.780 1.770 211.100 2.700 ;
        RECT 212.820 1.770 230.140 2.700 ;
        RECT 231.860 1.770 249.180 2.700 ;
        RECT 250.900 1.770 268.220 2.700 ;
        RECT 269.940 1.770 287.260 2.700 ;
        RECT 288.980 1.770 306.300 2.700 ;
        RECT 308.020 1.770 325.340 2.700 ;
        RECT 327.060 1.770 344.380 2.700 ;
        RECT 346.100 1.770 363.420 2.700 ;
        RECT 365.140 1.770 382.460 2.700 ;
        RECT 384.180 1.770 401.500 2.700 ;
        RECT 403.220 1.770 420.540 2.700 ;
        RECT 422.260 1.770 439.580 2.700 ;
        RECT 441.300 1.770 458.620 2.700 ;
        RECT 460.340 1.770 477.660 2.700 ;
        RECT 479.380 1.770 496.700 2.700 ;
        RECT 498.420 1.770 515.740 2.700 ;
        RECT 517.460 1.770 534.780 2.700 ;
        RECT 536.500 1.770 553.820 2.700 ;
        RECT 555.540 1.770 572.860 2.700 ;
        RECT 574.580 1.770 591.900 2.700 ;
        RECT 593.620 1.770 610.940 2.700 ;
        RECT 612.660 1.770 629.980 2.700 ;
        RECT 631.700 1.770 649.020 2.700 ;
        RECT 650.740 1.770 668.060 2.700 ;
        RECT 669.780 1.770 687.100 2.700 ;
        RECT 688.820 1.770 706.140 2.700 ;
        RECT 707.860 1.770 725.180 2.700 ;
        RECT 726.900 1.770 744.220 2.700 ;
        RECT 745.940 1.770 763.260 2.700 ;
        RECT 764.980 1.770 782.300 2.700 ;
        RECT 784.020 1.770 801.340 2.700 ;
        RECT 803.060 1.770 820.380 2.700 ;
        RECT 822.100 1.770 839.420 2.700 ;
        RECT 841.140 1.770 858.460 2.700 ;
        RECT 860.180 1.770 877.500 2.700 ;
        RECT 879.220 1.770 891.940 2.700 ;
      LAYER Metal3 ;
        RECT 9.610 1.820 891.990 701.820 ;
      LAYER Metal4 ;
        RECT 32.620 15.080 189.870 659.590 ;
        RECT 193.570 15.080 208.470 659.590 ;
        RECT 212.170 15.080 369.870 659.590 ;
        RECT 373.570 15.080 388.470 659.590 ;
        RECT 392.170 15.080 549.870 659.590 ;
        RECT 553.570 15.080 568.470 659.590 ;
        RECT 572.170 15.080 729.870 659.590 ;
        RECT 733.570 15.080 748.470 659.590 ;
        RECT 752.170 15.080 865.620 659.590 ;
        RECT 32.620 4.570 865.620 15.080 ;
  END
END driver_core
END LIBRARY

