magic
tech gf180mcuC
magscale 1 5
timestamp 1670065060
<< obsm1 >>
rect 672 1538 24304 23158
<< metal2 >>
rect 6188 -480 6300 240
rect 18676 -480 18788 240
<< obsm2 >>
rect 910 270 22274 23147
rect 910 196 6158 270
rect 6330 196 18646 270
rect 18818 196 22274 270
<< metal3 >>
rect -480 20692 240 20804
rect -480 12404 240 12516
rect 24760 12404 25480 12516
rect -480 4116 240 4228
<< obsm3 >>
rect 196 20834 24760 23142
rect 270 20662 24760 20834
rect 196 12546 24760 20662
rect 270 12374 24730 12546
rect 196 4258 24760 12374
rect 270 4086 24760 4258
rect 196 1554 24760 4086
<< metal4 >>
rect 1017 1538 1327 23158
rect 2877 1538 3187 23158
rect 19017 1538 19327 23158
rect 20877 1538 21187 23158
<< labels >>
rlabel metal3 s -480 4116 240 4228 4 clock_out_a
port 1 nsew signal output
rlabel metal3 s -480 12404 240 12516 4 clock_out_b
port 2 nsew signal output
rlabel metal3 s -480 20692 240 20804 4 clock_out_c
port 3 nsew signal output
rlabel metal2 s 6188 -480 6300 240 8 core_clock
port 4 nsew signal input
rlabel metal3 s 24760 12404 25480 12516 6 io_clock
port 5 nsew signal input
rlabel metal2 s 18676 -480 18788 240 8 la_oenb
port 6 nsew signal input
rlabel metal4 s 1017 1538 1327 23158 6 vccd1
port 7 nsew power bidirectional
rlabel metal4 s 19017 1538 19327 23158 6 vccd1
port 7 nsew power bidirectional
rlabel metal4 s 2877 1538 3187 23158 6 vssd1
port 8 nsew ground bidirectional
rlabel metal4 s 20877 1538 21187 23158 6 vssd1
port 8 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 25000 25000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 373392
string GDS_FILE /home/jasteve4/Documents/MicroMotorSequencerGL180/openlane/clock_source_sel/runs/22_12_03_05_56/results/signoff/clock_source_sel.magic.gds
string GDS_START 77534
<< end >>

