magic
tech gf180mcuC
magscale 1 5
timestamp 1670065060
<< metal1 >>
rect 672 23141 24304 23158
rect 672 23115 1029 23141
rect 1055 23115 1081 23141
rect 1107 23115 1133 23141
rect 1159 23115 1185 23141
rect 1211 23115 1237 23141
rect 1263 23115 1289 23141
rect 1315 23115 19029 23141
rect 19055 23115 19081 23141
rect 19107 23115 19133 23141
rect 19159 23115 19185 23141
rect 19211 23115 19237 23141
rect 19263 23115 19289 23141
rect 19315 23115 24304 23141
rect 672 23098 24304 23115
rect 672 22749 24304 22766
rect 672 22723 2889 22749
rect 2915 22723 2941 22749
rect 2967 22723 2993 22749
rect 3019 22723 3045 22749
rect 3071 22723 3097 22749
rect 3123 22723 3149 22749
rect 3175 22723 20889 22749
rect 20915 22723 20941 22749
rect 20967 22723 20993 22749
rect 21019 22723 21045 22749
rect 21071 22723 21097 22749
rect 21123 22723 21149 22749
rect 21175 22723 24304 22749
rect 672 22706 24304 22723
rect 672 22357 24304 22374
rect 672 22331 1029 22357
rect 1055 22331 1081 22357
rect 1107 22331 1133 22357
rect 1159 22331 1185 22357
rect 1211 22331 1237 22357
rect 1263 22331 1289 22357
rect 1315 22331 19029 22357
rect 19055 22331 19081 22357
rect 19107 22331 19133 22357
rect 19159 22331 19185 22357
rect 19211 22331 19237 22357
rect 19263 22331 19289 22357
rect 19315 22331 24304 22357
rect 672 22314 24304 22331
rect 672 21965 24304 21982
rect 672 21939 2889 21965
rect 2915 21939 2941 21965
rect 2967 21939 2993 21965
rect 3019 21939 3045 21965
rect 3071 21939 3097 21965
rect 3123 21939 3149 21965
rect 3175 21939 20889 21965
rect 20915 21939 20941 21965
rect 20967 21939 20993 21965
rect 21019 21939 21045 21965
rect 21071 21939 21097 21965
rect 21123 21939 21149 21965
rect 21175 21939 24304 21965
rect 672 21922 24304 21939
rect 672 21573 24304 21590
rect 672 21547 1029 21573
rect 1055 21547 1081 21573
rect 1107 21547 1133 21573
rect 1159 21547 1185 21573
rect 1211 21547 1237 21573
rect 1263 21547 1289 21573
rect 1315 21547 19029 21573
rect 19055 21547 19081 21573
rect 19107 21547 19133 21573
rect 19159 21547 19185 21573
rect 19211 21547 19237 21573
rect 19263 21547 19289 21573
rect 19315 21547 24304 21573
rect 672 21530 24304 21547
rect 672 21181 24304 21198
rect 672 21155 2889 21181
rect 2915 21155 2941 21181
rect 2967 21155 2993 21181
rect 3019 21155 3045 21181
rect 3071 21155 3097 21181
rect 3123 21155 3149 21181
rect 3175 21155 20889 21181
rect 20915 21155 20941 21181
rect 20967 21155 20993 21181
rect 21019 21155 21045 21181
rect 21071 21155 21097 21181
rect 21123 21155 21149 21181
rect 21175 21155 24304 21181
rect 672 21138 24304 21155
rect 911 21041 937 21047
rect 911 21009 937 21015
rect 672 20789 24304 20806
rect 672 20763 1029 20789
rect 1055 20763 1081 20789
rect 1107 20763 1133 20789
rect 1159 20763 1185 20789
rect 1211 20763 1237 20789
rect 1263 20763 1289 20789
rect 1315 20763 19029 20789
rect 19055 20763 19081 20789
rect 19107 20763 19133 20789
rect 19159 20763 19185 20789
rect 19211 20763 19237 20789
rect 19263 20763 19289 20789
rect 19315 20763 24304 20789
rect 672 20746 24304 20763
rect 672 20397 24304 20414
rect 672 20371 2889 20397
rect 2915 20371 2941 20397
rect 2967 20371 2993 20397
rect 3019 20371 3045 20397
rect 3071 20371 3097 20397
rect 3123 20371 3149 20397
rect 3175 20371 20889 20397
rect 20915 20371 20941 20397
rect 20967 20371 20993 20397
rect 21019 20371 21045 20397
rect 21071 20371 21097 20397
rect 21123 20371 21149 20397
rect 21175 20371 24304 20397
rect 672 20354 24304 20371
rect 672 20005 24304 20022
rect 672 19979 1029 20005
rect 1055 19979 1081 20005
rect 1107 19979 1133 20005
rect 1159 19979 1185 20005
rect 1211 19979 1237 20005
rect 1263 19979 1289 20005
rect 1315 19979 19029 20005
rect 19055 19979 19081 20005
rect 19107 19979 19133 20005
rect 19159 19979 19185 20005
rect 19211 19979 19237 20005
rect 19263 19979 19289 20005
rect 19315 19979 24304 20005
rect 672 19962 24304 19979
rect 672 19613 24304 19630
rect 672 19587 2889 19613
rect 2915 19587 2941 19613
rect 2967 19587 2993 19613
rect 3019 19587 3045 19613
rect 3071 19587 3097 19613
rect 3123 19587 3149 19613
rect 3175 19587 20889 19613
rect 20915 19587 20941 19613
rect 20967 19587 20993 19613
rect 21019 19587 21045 19613
rect 21071 19587 21097 19613
rect 21123 19587 21149 19613
rect 21175 19587 24304 19613
rect 672 19570 24304 19587
rect 672 19221 24304 19238
rect 672 19195 1029 19221
rect 1055 19195 1081 19221
rect 1107 19195 1133 19221
rect 1159 19195 1185 19221
rect 1211 19195 1237 19221
rect 1263 19195 1289 19221
rect 1315 19195 19029 19221
rect 19055 19195 19081 19221
rect 19107 19195 19133 19221
rect 19159 19195 19185 19221
rect 19211 19195 19237 19221
rect 19263 19195 19289 19221
rect 19315 19195 24304 19221
rect 672 19178 24304 19195
rect 672 18829 24304 18846
rect 672 18803 2889 18829
rect 2915 18803 2941 18829
rect 2967 18803 2993 18829
rect 3019 18803 3045 18829
rect 3071 18803 3097 18829
rect 3123 18803 3149 18829
rect 3175 18803 20889 18829
rect 20915 18803 20941 18829
rect 20967 18803 20993 18829
rect 21019 18803 21045 18829
rect 21071 18803 21097 18829
rect 21123 18803 21149 18829
rect 21175 18803 24304 18829
rect 672 18786 24304 18803
rect 672 18437 24304 18454
rect 672 18411 1029 18437
rect 1055 18411 1081 18437
rect 1107 18411 1133 18437
rect 1159 18411 1185 18437
rect 1211 18411 1237 18437
rect 1263 18411 1289 18437
rect 1315 18411 19029 18437
rect 19055 18411 19081 18437
rect 19107 18411 19133 18437
rect 19159 18411 19185 18437
rect 19211 18411 19237 18437
rect 19263 18411 19289 18437
rect 19315 18411 24304 18437
rect 672 18394 24304 18411
rect 672 18045 24304 18062
rect 672 18019 2889 18045
rect 2915 18019 2941 18045
rect 2967 18019 2993 18045
rect 3019 18019 3045 18045
rect 3071 18019 3097 18045
rect 3123 18019 3149 18045
rect 3175 18019 20889 18045
rect 20915 18019 20941 18045
rect 20967 18019 20993 18045
rect 21019 18019 21045 18045
rect 21071 18019 21097 18045
rect 21123 18019 21149 18045
rect 21175 18019 24304 18045
rect 672 18002 24304 18019
rect 672 17653 24304 17670
rect 672 17627 1029 17653
rect 1055 17627 1081 17653
rect 1107 17627 1133 17653
rect 1159 17627 1185 17653
rect 1211 17627 1237 17653
rect 1263 17627 1289 17653
rect 1315 17627 19029 17653
rect 19055 17627 19081 17653
rect 19107 17627 19133 17653
rect 19159 17627 19185 17653
rect 19211 17627 19237 17653
rect 19263 17627 19289 17653
rect 19315 17627 24304 17653
rect 672 17610 24304 17627
rect 672 17261 24304 17278
rect 672 17235 2889 17261
rect 2915 17235 2941 17261
rect 2967 17235 2993 17261
rect 3019 17235 3045 17261
rect 3071 17235 3097 17261
rect 3123 17235 3149 17261
rect 3175 17235 20889 17261
rect 20915 17235 20941 17261
rect 20967 17235 20993 17261
rect 21019 17235 21045 17261
rect 21071 17235 21097 17261
rect 21123 17235 21149 17261
rect 21175 17235 24304 17261
rect 672 17218 24304 17235
rect 672 16869 24304 16886
rect 672 16843 1029 16869
rect 1055 16843 1081 16869
rect 1107 16843 1133 16869
rect 1159 16843 1185 16869
rect 1211 16843 1237 16869
rect 1263 16843 1289 16869
rect 1315 16843 19029 16869
rect 19055 16843 19081 16869
rect 19107 16843 19133 16869
rect 19159 16843 19185 16869
rect 19211 16843 19237 16869
rect 19263 16843 19289 16869
rect 19315 16843 24304 16869
rect 672 16826 24304 16843
rect 672 16477 24304 16494
rect 672 16451 2889 16477
rect 2915 16451 2941 16477
rect 2967 16451 2993 16477
rect 3019 16451 3045 16477
rect 3071 16451 3097 16477
rect 3123 16451 3149 16477
rect 3175 16451 20889 16477
rect 20915 16451 20941 16477
rect 20967 16451 20993 16477
rect 21019 16451 21045 16477
rect 21071 16451 21097 16477
rect 21123 16451 21149 16477
rect 21175 16451 24304 16477
rect 672 16434 24304 16451
rect 672 16085 24304 16102
rect 672 16059 1029 16085
rect 1055 16059 1081 16085
rect 1107 16059 1133 16085
rect 1159 16059 1185 16085
rect 1211 16059 1237 16085
rect 1263 16059 1289 16085
rect 1315 16059 19029 16085
rect 19055 16059 19081 16085
rect 19107 16059 19133 16085
rect 19159 16059 19185 16085
rect 19211 16059 19237 16085
rect 19263 16059 19289 16085
rect 19315 16059 24304 16085
rect 672 16042 24304 16059
rect 672 15693 24304 15710
rect 672 15667 2889 15693
rect 2915 15667 2941 15693
rect 2967 15667 2993 15693
rect 3019 15667 3045 15693
rect 3071 15667 3097 15693
rect 3123 15667 3149 15693
rect 3175 15667 20889 15693
rect 20915 15667 20941 15693
rect 20967 15667 20993 15693
rect 21019 15667 21045 15693
rect 21071 15667 21097 15693
rect 21123 15667 21149 15693
rect 21175 15667 24304 15693
rect 672 15650 24304 15667
rect 672 15301 24304 15318
rect 672 15275 1029 15301
rect 1055 15275 1081 15301
rect 1107 15275 1133 15301
rect 1159 15275 1185 15301
rect 1211 15275 1237 15301
rect 1263 15275 1289 15301
rect 1315 15275 19029 15301
rect 19055 15275 19081 15301
rect 19107 15275 19133 15301
rect 19159 15275 19185 15301
rect 19211 15275 19237 15301
rect 19263 15275 19289 15301
rect 19315 15275 24304 15301
rect 672 15258 24304 15275
rect 672 14909 24304 14926
rect 672 14883 2889 14909
rect 2915 14883 2941 14909
rect 2967 14883 2993 14909
rect 3019 14883 3045 14909
rect 3071 14883 3097 14909
rect 3123 14883 3149 14909
rect 3175 14883 20889 14909
rect 20915 14883 20941 14909
rect 20967 14883 20993 14909
rect 21019 14883 21045 14909
rect 21071 14883 21097 14909
rect 21123 14883 21149 14909
rect 21175 14883 24304 14909
rect 672 14866 24304 14883
rect 672 14517 24304 14534
rect 672 14491 1029 14517
rect 1055 14491 1081 14517
rect 1107 14491 1133 14517
rect 1159 14491 1185 14517
rect 1211 14491 1237 14517
rect 1263 14491 1289 14517
rect 1315 14491 19029 14517
rect 19055 14491 19081 14517
rect 19107 14491 19133 14517
rect 19159 14491 19185 14517
rect 19211 14491 19237 14517
rect 19263 14491 19289 14517
rect 19315 14491 24304 14517
rect 672 14474 24304 14491
rect 672 14125 24304 14142
rect 672 14099 2889 14125
rect 2915 14099 2941 14125
rect 2967 14099 2993 14125
rect 3019 14099 3045 14125
rect 3071 14099 3097 14125
rect 3123 14099 3149 14125
rect 3175 14099 20889 14125
rect 20915 14099 20941 14125
rect 20967 14099 20993 14125
rect 21019 14099 21045 14125
rect 21071 14099 21097 14125
rect 21123 14099 21149 14125
rect 21175 14099 24304 14125
rect 672 14082 24304 14099
rect 672 13733 24304 13750
rect 672 13707 1029 13733
rect 1055 13707 1081 13733
rect 1107 13707 1133 13733
rect 1159 13707 1185 13733
rect 1211 13707 1237 13733
rect 1263 13707 1289 13733
rect 1315 13707 19029 13733
rect 19055 13707 19081 13733
rect 19107 13707 19133 13733
rect 19159 13707 19185 13733
rect 19211 13707 19237 13733
rect 19263 13707 19289 13733
rect 19315 13707 24304 13733
rect 672 13690 24304 13707
rect 672 13341 24304 13358
rect 672 13315 2889 13341
rect 2915 13315 2941 13341
rect 2967 13315 2993 13341
rect 3019 13315 3045 13341
rect 3071 13315 3097 13341
rect 3123 13315 3149 13341
rect 3175 13315 20889 13341
rect 20915 13315 20941 13341
rect 20967 13315 20993 13341
rect 21019 13315 21045 13341
rect 21071 13315 21097 13341
rect 21123 13315 21149 13341
rect 21175 13315 24304 13341
rect 672 13298 24304 13315
rect 672 12949 24304 12966
rect 672 12923 1029 12949
rect 1055 12923 1081 12949
rect 1107 12923 1133 12949
rect 1159 12923 1185 12949
rect 1211 12923 1237 12949
rect 1263 12923 1289 12949
rect 1315 12923 19029 12949
rect 19055 12923 19081 12949
rect 19107 12923 19133 12949
rect 19159 12923 19185 12949
rect 19211 12923 19237 12949
rect 19263 12923 19289 12949
rect 19315 12923 24304 12949
rect 672 12906 24304 12923
rect 911 12641 937 12647
rect 911 12609 937 12615
rect 672 12557 24304 12574
rect 672 12531 2889 12557
rect 2915 12531 2941 12557
rect 2967 12531 2993 12557
rect 3019 12531 3045 12557
rect 3071 12531 3097 12557
rect 3123 12531 3149 12557
rect 3175 12531 20889 12557
rect 20915 12531 20941 12557
rect 20967 12531 20993 12557
rect 21019 12531 21045 12557
rect 21071 12531 21097 12557
rect 21123 12531 21149 12557
rect 21175 12531 24304 12557
rect 672 12514 24304 12531
rect 672 12165 24304 12182
rect 672 12139 1029 12165
rect 1055 12139 1081 12165
rect 1107 12139 1133 12165
rect 1159 12139 1185 12165
rect 1211 12139 1237 12165
rect 1263 12139 1289 12165
rect 1315 12139 19029 12165
rect 19055 12139 19081 12165
rect 19107 12139 19133 12165
rect 19159 12139 19185 12165
rect 19211 12139 19237 12165
rect 19263 12139 19289 12165
rect 19315 12139 24304 12165
rect 672 12122 24304 12139
rect 672 11773 24304 11790
rect 672 11747 2889 11773
rect 2915 11747 2941 11773
rect 2967 11747 2993 11773
rect 3019 11747 3045 11773
rect 3071 11747 3097 11773
rect 3123 11747 3149 11773
rect 3175 11747 20889 11773
rect 20915 11747 20941 11773
rect 20967 11747 20993 11773
rect 21019 11747 21045 11773
rect 21071 11747 21097 11773
rect 21123 11747 21149 11773
rect 21175 11747 24304 11773
rect 672 11730 24304 11747
rect 672 11381 24304 11398
rect 672 11355 1029 11381
rect 1055 11355 1081 11381
rect 1107 11355 1133 11381
rect 1159 11355 1185 11381
rect 1211 11355 1237 11381
rect 1263 11355 1289 11381
rect 1315 11355 19029 11381
rect 19055 11355 19081 11381
rect 19107 11355 19133 11381
rect 19159 11355 19185 11381
rect 19211 11355 19237 11381
rect 19263 11355 19289 11381
rect 19315 11355 24304 11381
rect 672 11338 24304 11355
rect 672 10989 24304 11006
rect 672 10963 2889 10989
rect 2915 10963 2941 10989
rect 2967 10963 2993 10989
rect 3019 10963 3045 10989
rect 3071 10963 3097 10989
rect 3123 10963 3149 10989
rect 3175 10963 20889 10989
rect 20915 10963 20941 10989
rect 20967 10963 20993 10989
rect 21019 10963 21045 10989
rect 21071 10963 21097 10989
rect 21123 10963 21149 10989
rect 21175 10963 24304 10989
rect 672 10946 24304 10963
rect 672 10597 24304 10614
rect 672 10571 1029 10597
rect 1055 10571 1081 10597
rect 1107 10571 1133 10597
rect 1159 10571 1185 10597
rect 1211 10571 1237 10597
rect 1263 10571 1289 10597
rect 1315 10571 19029 10597
rect 19055 10571 19081 10597
rect 19107 10571 19133 10597
rect 19159 10571 19185 10597
rect 19211 10571 19237 10597
rect 19263 10571 19289 10597
rect 19315 10571 24304 10597
rect 672 10554 24304 10571
rect 672 10205 24304 10222
rect 672 10179 2889 10205
rect 2915 10179 2941 10205
rect 2967 10179 2993 10205
rect 3019 10179 3045 10205
rect 3071 10179 3097 10205
rect 3123 10179 3149 10205
rect 3175 10179 20889 10205
rect 20915 10179 20941 10205
rect 20967 10179 20993 10205
rect 21019 10179 21045 10205
rect 21071 10179 21097 10205
rect 21123 10179 21149 10205
rect 21175 10179 24304 10205
rect 672 10162 24304 10179
rect 672 9813 24304 9830
rect 672 9787 1029 9813
rect 1055 9787 1081 9813
rect 1107 9787 1133 9813
rect 1159 9787 1185 9813
rect 1211 9787 1237 9813
rect 1263 9787 1289 9813
rect 1315 9787 19029 9813
rect 19055 9787 19081 9813
rect 19107 9787 19133 9813
rect 19159 9787 19185 9813
rect 19211 9787 19237 9813
rect 19263 9787 19289 9813
rect 19315 9787 24304 9813
rect 672 9770 24304 9787
rect 672 9421 24304 9438
rect 672 9395 2889 9421
rect 2915 9395 2941 9421
rect 2967 9395 2993 9421
rect 3019 9395 3045 9421
rect 3071 9395 3097 9421
rect 3123 9395 3149 9421
rect 3175 9395 20889 9421
rect 20915 9395 20941 9421
rect 20967 9395 20993 9421
rect 21019 9395 21045 9421
rect 21071 9395 21097 9421
rect 21123 9395 21149 9421
rect 21175 9395 24304 9421
rect 672 9378 24304 9395
rect 672 9029 24304 9046
rect 672 9003 1029 9029
rect 1055 9003 1081 9029
rect 1107 9003 1133 9029
rect 1159 9003 1185 9029
rect 1211 9003 1237 9029
rect 1263 9003 1289 9029
rect 1315 9003 19029 9029
rect 19055 9003 19081 9029
rect 19107 9003 19133 9029
rect 19159 9003 19185 9029
rect 19211 9003 19237 9029
rect 19263 9003 19289 9029
rect 19315 9003 24304 9029
rect 672 8986 24304 9003
rect 672 8637 24304 8654
rect 672 8611 2889 8637
rect 2915 8611 2941 8637
rect 2967 8611 2993 8637
rect 3019 8611 3045 8637
rect 3071 8611 3097 8637
rect 3123 8611 3149 8637
rect 3175 8611 20889 8637
rect 20915 8611 20941 8637
rect 20967 8611 20993 8637
rect 21019 8611 21045 8637
rect 21071 8611 21097 8637
rect 21123 8611 21149 8637
rect 21175 8611 24304 8637
rect 672 8594 24304 8611
rect 672 8245 24304 8262
rect 672 8219 1029 8245
rect 1055 8219 1081 8245
rect 1107 8219 1133 8245
rect 1159 8219 1185 8245
rect 1211 8219 1237 8245
rect 1263 8219 1289 8245
rect 1315 8219 19029 8245
rect 19055 8219 19081 8245
rect 19107 8219 19133 8245
rect 19159 8219 19185 8245
rect 19211 8219 19237 8245
rect 19263 8219 19289 8245
rect 19315 8219 24304 8245
rect 672 8202 24304 8219
rect 672 7853 24304 7870
rect 672 7827 2889 7853
rect 2915 7827 2941 7853
rect 2967 7827 2993 7853
rect 3019 7827 3045 7853
rect 3071 7827 3097 7853
rect 3123 7827 3149 7853
rect 3175 7827 20889 7853
rect 20915 7827 20941 7853
rect 20967 7827 20993 7853
rect 21019 7827 21045 7853
rect 21071 7827 21097 7853
rect 21123 7827 21149 7853
rect 21175 7827 24304 7853
rect 672 7810 24304 7827
rect 672 7461 24304 7478
rect 672 7435 1029 7461
rect 1055 7435 1081 7461
rect 1107 7435 1133 7461
rect 1159 7435 1185 7461
rect 1211 7435 1237 7461
rect 1263 7435 1289 7461
rect 1315 7435 19029 7461
rect 19055 7435 19081 7461
rect 19107 7435 19133 7461
rect 19159 7435 19185 7461
rect 19211 7435 19237 7461
rect 19263 7435 19289 7461
rect 19315 7435 24304 7461
rect 672 7418 24304 7435
rect 672 7069 24304 7086
rect 672 7043 2889 7069
rect 2915 7043 2941 7069
rect 2967 7043 2993 7069
rect 3019 7043 3045 7069
rect 3071 7043 3097 7069
rect 3123 7043 3149 7069
rect 3175 7043 20889 7069
rect 20915 7043 20941 7069
rect 20967 7043 20993 7069
rect 21019 7043 21045 7069
rect 21071 7043 21097 7069
rect 21123 7043 21149 7069
rect 21175 7043 24304 7069
rect 672 7026 24304 7043
rect 672 6677 24304 6694
rect 672 6651 1029 6677
rect 1055 6651 1081 6677
rect 1107 6651 1133 6677
rect 1159 6651 1185 6677
rect 1211 6651 1237 6677
rect 1263 6651 1289 6677
rect 1315 6651 19029 6677
rect 19055 6651 19081 6677
rect 19107 6651 19133 6677
rect 19159 6651 19185 6677
rect 19211 6651 19237 6677
rect 19263 6651 19289 6677
rect 19315 6651 24304 6677
rect 672 6634 24304 6651
rect 672 6285 24304 6302
rect 672 6259 2889 6285
rect 2915 6259 2941 6285
rect 2967 6259 2993 6285
rect 3019 6259 3045 6285
rect 3071 6259 3097 6285
rect 3123 6259 3149 6285
rect 3175 6259 20889 6285
rect 20915 6259 20941 6285
rect 20967 6259 20993 6285
rect 21019 6259 21045 6285
rect 21071 6259 21097 6285
rect 21123 6259 21149 6285
rect 21175 6259 24304 6285
rect 672 6242 24304 6259
rect 16255 6089 16281 6095
rect 16025 6063 16031 6089
rect 16057 6063 16063 6089
rect 16255 6057 16281 6063
rect 13505 6007 13511 6033
rect 13537 6007 13543 6033
rect 672 5893 24304 5910
rect 672 5867 1029 5893
rect 1055 5867 1081 5893
rect 1107 5867 1133 5893
rect 1159 5867 1185 5893
rect 1211 5867 1237 5893
rect 1263 5867 1289 5893
rect 1315 5867 19029 5893
rect 19055 5867 19081 5893
rect 19107 5867 19133 5893
rect 19159 5867 19185 5893
rect 19211 5867 19237 5893
rect 19263 5867 19289 5893
rect 19315 5867 24304 5893
rect 672 5850 24304 5867
rect 12503 5697 12529 5703
rect 12833 5671 12839 5697
rect 12865 5671 12871 5697
rect 12503 5665 12529 5671
rect 12889 5615 12895 5641
rect 12921 5615 12927 5641
rect 12335 5585 12361 5591
rect 12335 5553 12361 5559
rect 13231 5585 13257 5591
rect 13231 5553 13257 5559
rect 672 5501 24304 5518
rect 672 5475 2889 5501
rect 2915 5475 2941 5501
rect 2967 5475 2993 5501
rect 3019 5475 3045 5501
rect 3071 5475 3097 5501
rect 3123 5475 3149 5501
rect 3175 5475 20889 5501
rect 20915 5475 20941 5501
rect 20967 5475 20993 5501
rect 21019 5475 21045 5501
rect 21071 5475 21097 5501
rect 21123 5475 21149 5501
rect 21175 5475 24304 5501
rect 672 5458 24304 5475
rect 11887 5417 11913 5423
rect 11887 5385 11913 5391
rect 11713 5335 11719 5361
rect 11745 5335 11751 5361
rect 12833 5279 12839 5305
rect 12865 5279 12871 5305
rect 12503 5249 12529 5255
rect 14289 5223 14295 5249
rect 14321 5223 14327 5249
rect 12503 5217 12529 5223
rect 672 5109 24304 5126
rect 672 5083 1029 5109
rect 1055 5083 1081 5109
rect 1107 5083 1133 5109
rect 1159 5083 1185 5109
rect 1211 5083 1237 5109
rect 1263 5083 1289 5109
rect 1315 5083 19029 5109
rect 19055 5083 19081 5109
rect 19107 5083 19133 5109
rect 19159 5083 19185 5109
rect 19211 5083 19237 5109
rect 19263 5083 19289 5109
rect 19315 5083 24304 5109
rect 672 5066 24304 5083
rect 13337 4943 13343 4969
rect 13369 4943 13375 4969
rect 11881 4887 11887 4913
rect 11913 4887 11919 4913
rect 12273 4831 12279 4857
rect 12305 4831 12311 4857
rect 13567 4801 13593 4807
rect 13567 4769 13593 4775
rect 672 4717 24304 4734
rect 672 4691 2889 4717
rect 2915 4691 2941 4717
rect 2967 4691 2993 4717
rect 3019 4691 3045 4717
rect 3071 4691 3097 4717
rect 3123 4691 3149 4717
rect 3175 4691 20889 4717
rect 20915 4691 20941 4717
rect 20967 4691 20993 4717
rect 21019 4691 21045 4717
rect 21071 4691 21097 4717
rect 21123 4691 21149 4717
rect 21175 4691 24304 4717
rect 672 4674 24304 4691
rect 905 4551 911 4577
rect 937 4551 943 4577
rect 1079 4521 1105 4527
rect 1079 4489 1105 4495
rect 1359 4521 1385 4527
rect 1359 4489 1385 4495
rect 672 4325 24304 4342
rect 672 4299 1029 4325
rect 1055 4299 1081 4325
rect 1107 4299 1133 4325
rect 1159 4299 1185 4325
rect 1211 4299 1237 4325
rect 1263 4299 1289 4325
rect 1315 4299 19029 4325
rect 19055 4299 19081 4325
rect 19107 4299 19133 4325
rect 19159 4299 19185 4325
rect 19211 4299 19237 4325
rect 19263 4299 19289 4325
rect 19315 4299 24304 4325
rect 672 4282 24304 4299
rect 672 3933 24304 3950
rect 672 3907 2889 3933
rect 2915 3907 2941 3933
rect 2967 3907 2993 3933
rect 3019 3907 3045 3933
rect 3071 3907 3097 3933
rect 3123 3907 3149 3933
rect 3175 3907 20889 3933
rect 20915 3907 20941 3933
rect 20967 3907 20993 3933
rect 21019 3907 21045 3933
rect 21071 3907 21097 3933
rect 21123 3907 21149 3933
rect 21175 3907 24304 3933
rect 672 3890 24304 3907
rect 10873 3767 10879 3793
rect 10905 3767 10911 3793
rect 12447 3737 12473 3743
rect 12217 3711 12223 3737
rect 12249 3711 12255 3737
rect 12447 3705 12473 3711
rect 672 3541 24304 3558
rect 672 3515 1029 3541
rect 1055 3515 1081 3541
rect 1107 3515 1133 3541
rect 1159 3515 1185 3541
rect 1211 3515 1237 3541
rect 1263 3515 1289 3541
rect 1315 3515 19029 3541
rect 19055 3515 19081 3541
rect 19107 3515 19133 3541
rect 19159 3515 19185 3541
rect 19211 3515 19237 3541
rect 19263 3515 19289 3541
rect 19315 3515 24304 3541
rect 672 3498 24304 3515
rect 672 3149 24304 3166
rect 672 3123 2889 3149
rect 2915 3123 2941 3149
rect 2967 3123 2993 3149
rect 3019 3123 3045 3149
rect 3071 3123 3097 3149
rect 3123 3123 3149 3149
rect 3175 3123 20889 3149
rect 20915 3123 20941 3149
rect 20967 3123 20993 3149
rect 21019 3123 21045 3149
rect 21071 3123 21097 3149
rect 21123 3123 21149 3149
rect 21175 3123 24304 3149
rect 672 3106 24304 3123
rect 672 2757 24304 2774
rect 672 2731 1029 2757
rect 1055 2731 1081 2757
rect 1107 2731 1133 2757
rect 1159 2731 1185 2757
rect 1211 2731 1237 2757
rect 1263 2731 1289 2757
rect 1315 2731 19029 2757
rect 19055 2731 19081 2757
rect 19107 2731 19133 2757
rect 19159 2731 19185 2757
rect 19211 2731 19237 2757
rect 19263 2731 19289 2757
rect 19315 2731 24304 2757
rect 672 2714 24304 2731
rect 672 2365 24304 2382
rect 672 2339 2889 2365
rect 2915 2339 2941 2365
rect 2967 2339 2993 2365
rect 3019 2339 3045 2365
rect 3071 2339 3097 2365
rect 3123 2339 3149 2365
rect 3175 2339 20889 2365
rect 20915 2339 20941 2365
rect 20967 2339 20993 2365
rect 21019 2339 21045 2365
rect 21071 2339 21097 2365
rect 21123 2339 21149 2365
rect 21175 2339 24304 2365
rect 672 2322 24304 2339
rect 672 1973 24304 1990
rect 672 1947 1029 1973
rect 1055 1947 1081 1973
rect 1107 1947 1133 1973
rect 1159 1947 1185 1973
rect 1211 1947 1237 1973
rect 1263 1947 1289 1973
rect 1315 1947 19029 1973
rect 19055 1947 19081 1973
rect 19107 1947 19133 1973
rect 19159 1947 19185 1973
rect 19211 1947 19237 1973
rect 19263 1947 19289 1973
rect 19315 1947 24304 1973
rect 672 1930 24304 1947
rect 18607 1721 18633 1727
rect 18607 1689 18633 1695
rect 18999 1721 19025 1727
rect 18999 1689 19025 1695
rect 18831 1665 18857 1671
rect 18831 1633 18857 1639
rect 672 1581 24304 1598
rect 672 1555 2889 1581
rect 2915 1555 2941 1581
rect 2967 1555 2993 1581
rect 3019 1555 3045 1581
rect 3071 1555 3097 1581
rect 3123 1555 3149 1581
rect 3175 1555 20889 1581
rect 20915 1555 20941 1581
rect 20967 1555 20993 1581
rect 21019 1555 21045 1581
rect 21071 1555 21097 1581
rect 21123 1555 21149 1581
rect 21175 1555 24304 1581
rect 672 1538 24304 1555
<< via1 >>
rect 1029 23115 1055 23141
rect 1081 23115 1107 23141
rect 1133 23115 1159 23141
rect 1185 23115 1211 23141
rect 1237 23115 1263 23141
rect 1289 23115 1315 23141
rect 19029 23115 19055 23141
rect 19081 23115 19107 23141
rect 19133 23115 19159 23141
rect 19185 23115 19211 23141
rect 19237 23115 19263 23141
rect 19289 23115 19315 23141
rect 2889 22723 2915 22749
rect 2941 22723 2967 22749
rect 2993 22723 3019 22749
rect 3045 22723 3071 22749
rect 3097 22723 3123 22749
rect 3149 22723 3175 22749
rect 20889 22723 20915 22749
rect 20941 22723 20967 22749
rect 20993 22723 21019 22749
rect 21045 22723 21071 22749
rect 21097 22723 21123 22749
rect 21149 22723 21175 22749
rect 1029 22331 1055 22357
rect 1081 22331 1107 22357
rect 1133 22331 1159 22357
rect 1185 22331 1211 22357
rect 1237 22331 1263 22357
rect 1289 22331 1315 22357
rect 19029 22331 19055 22357
rect 19081 22331 19107 22357
rect 19133 22331 19159 22357
rect 19185 22331 19211 22357
rect 19237 22331 19263 22357
rect 19289 22331 19315 22357
rect 2889 21939 2915 21965
rect 2941 21939 2967 21965
rect 2993 21939 3019 21965
rect 3045 21939 3071 21965
rect 3097 21939 3123 21965
rect 3149 21939 3175 21965
rect 20889 21939 20915 21965
rect 20941 21939 20967 21965
rect 20993 21939 21019 21965
rect 21045 21939 21071 21965
rect 21097 21939 21123 21965
rect 21149 21939 21175 21965
rect 1029 21547 1055 21573
rect 1081 21547 1107 21573
rect 1133 21547 1159 21573
rect 1185 21547 1211 21573
rect 1237 21547 1263 21573
rect 1289 21547 1315 21573
rect 19029 21547 19055 21573
rect 19081 21547 19107 21573
rect 19133 21547 19159 21573
rect 19185 21547 19211 21573
rect 19237 21547 19263 21573
rect 19289 21547 19315 21573
rect 2889 21155 2915 21181
rect 2941 21155 2967 21181
rect 2993 21155 3019 21181
rect 3045 21155 3071 21181
rect 3097 21155 3123 21181
rect 3149 21155 3175 21181
rect 20889 21155 20915 21181
rect 20941 21155 20967 21181
rect 20993 21155 21019 21181
rect 21045 21155 21071 21181
rect 21097 21155 21123 21181
rect 21149 21155 21175 21181
rect 911 21015 937 21041
rect 1029 20763 1055 20789
rect 1081 20763 1107 20789
rect 1133 20763 1159 20789
rect 1185 20763 1211 20789
rect 1237 20763 1263 20789
rect 1289 20763 1315 20789
rect 19029 20763 19055 20789
rect 19081 20763 19107 20789
rect 19133 20763 19159 20789
rect 19185 20763 19211 20789
rect 19237 20763 19263 20789
rect 19289 20763 19315 20789
rect 2889 20371 2915 20397
rect 2941 20371 2967 20397
rect 2993 20371 3019 20397
rect 3045 20371 3071 20397
rect 3097 20371 3123 20397
rect 3149 20371 3175 20397
rect 20889 20371 20915 20397
rect 20941 20371 20967 20397
rect 20993 20371 21019 20397
rect 21045 20371 21071 20397
rect 21097 20371 21123 20397
rect 21149 20371 21175 20397
rect 1029 19979 1055 20005
rect 1081 19979 1107 20005
rect 1133 19979 1159 20005
rect 1185 19979 1211 20005
rect 1237 19979 1263 20005
rect 1289 19979 1315 20005
rect 19029 19979 19055 20005
rect 19081 19979 19107 20005
rect 19133 19979 19159 20005
rect 19185 19979 19211 20005
rect 19237 19979 19263 20005
rect 19289 19979 19315 20005
rect 2889 19587 2915 19613
rect 2941 19587 2967 19613
rect 2993 19587 3019 19613
rect 3045 19587 3071 19613
rect 3097 19587 3123 19613
rect 3149 19587 3175 19613
rect 20889 19587 20915 19613
rect 20941 19587 20967 19613
rect 20993 19587 21019 19613
rect 21045 19587 21071 19613
rect 21097 19587 21123 19613
rect 21149 19587 21175 19613
rect 1029 19195 1055 19221
rect 1081 19195 1107 19221
rect 1133 19195 1159 19221
rect 1185 19195 1211 19221
rect 1237 19195 1263 19221
rect 1289 19195 1315 19221
rect 19029 19195 19055 19221
rect 19081 19195 19107 19221
rect 19133 19195 19159 19221
rect 19185 19195 19211 19221
rect 19237 19195 19263 19221
rect 19289 19195 19315 19221
rect 2889 18803 2915 18829
rect 2941 18803 2967 18829
rect 2993 18803 3019 18829
rect 3045 18803 3071 18829
rect 3097 18803 3123 18829
rect 3149 18803 3175 18829
rect 20889 18803 20915 18829
rect 20941 18803 20967 18829
rect 20993 18803 21019 18829
rect 21045 18803 21071 18829
rect 21097 18803 21123 18829
rect 21149 18803 21175 18829
rect 1029 18411 1055 18437
rect 1081 18411 1107 18437
rect 1133 18411 1159 18437
rect 1185 18411 1211 18437
rect 1237 18411 1263 18437
rect 1289 18411 1315 18437
rect 19029 18411 19055 18437
rect 19081 18411 19107 18437
rect 19133 18411 19159 18437
rect 19185 18411 19211 18437
rect 19237 18411 19263 18437
rect 19289 18411 19315 18437
rect 2889 18019 2915 18045
rect 2941 18019 2967 18045
rect 2993 18019 3019 18045
rect 3045 18019 3071 18045
rect 3097 18019 3123 18045
rect 3149 18019 3175 18045
rect 20889 18019 20915 18045
rect 20941 18019 20967 18045
rect 20993 18019 21019 18045
rect 21045 18019 21071 18045
rect 21097 18019 21123 18045
rect 21149 18019 21175 18045
rect 1029 17627 1055 17653
rect 1081 17627 1107 17653
rect 1133 17627 1159 17653
rect 1185 17627 1211 17653
rect 1237 17627 1263 17653
rect 1289 17627 1315 17653
rect 19029 17627 19055 17653
rect 19081 17627 19107 17653
rect 19133 17627 19159 17653
rect 19185 17627 19211 17653
rect 19237 17627 19263 17653
rect 19289 17627 19315 17653
rect 2889 17235 2915 17261
rect 2941 17235 2967 17261
rect 2993 17235 3019 17261
rect 3045 17235 3071 17261
rect 3097 17235 3123 17261
rect 3149 17235 3175 17261
rect 20889 17235 20915 17261
rect 20941 17235 20967 17261
rect 20993 17235 21019 17261
rect 21045 17235 21071 17261
rect 21097 17235 21123 17261
rect 21149 17235 21175 17261
rect 1029 16843 1055 16869
rect 1081 16843 1107 16869
rect 1133 16843 1159 16869
rect 1185 16843 1211 16869
rect 1237 16843 1263 16869
rect 1289 16843 1315 16869
rect 19029 16843 19055 16869
rect 19081 16843 19107 16869
rect 19133 16843 19159 16869
rect 19185 16843 19211 16869
rect 19237 16843 19263 16869
rect 19289 16843 19315 16869
rect 2889 16451 2915 16477
rect 2941 16451 2967 16477
rect 2993 16451 3019 16477
rect 3045 16451 3071 16477
rect 3097 16451 3123 16477
rect 3149 16451 3175 16477
rect 20889 16451 20915 16477
rect 20941 16451 20967 16477
rect 20993 16451 21019 16477
rect 21045 16451 21071 16477
rect 21097 16451 21123 16477
rect 21149 16451 21175 16477
rect 1029 16059 1055 16085
rect 1081 16059 1107 16085
rect 1133 16059 1159 16085
rect 1185 16059 1211 16085
rect 1237 16059 1263 16085
rect 1289 16059 1315 16085
rect 19029 16059 19055 16085
rect 19081 16059 19107 16085
rect 19133 16059 19159 16085
rect 19185 16059 19211 16085
rect 19237 16059 19263 16085
rect 19289 16059 19315 16085
rect 2889 15667 2915 15693
rect 2941 15667 2967 15693
rect 2993 15667 3019 15693
rect 3045 15667 3071 15693
rect 3097 15667 3123 15693
rect 3149 15667 3175 15693
rect 20889 15667 20915 15693
rect 20941 15667 20967 15693
rect 20993 15667 21019 15693
rect 21045 15667 21071 15693
rect 21097 15667 21123 15693
rect 21149 15667 21175 15693
rect 1029 15275 1055 15301
rect 1081 15275 1107 15301
rect 1133 15275 1159 15301
rect 1185 15275 1211 15301
rect 1237 15275 1263 15301
rect 1289 15275 1315 15301
rect 19029 15275 19055 15301
rect 19081 15275 19107 15301
rect 19133 15275 19159 15301
rect 19185 15275 19211 15301
rect 19237 15275 19263 15301
rect 19289 15275 19315 15301
rect 2889 14883 2915 14909
rect 2941 14883 2967 14909
rect 2993 14883 3019 14909
rect 3045 14883 3071 14909
rect 3097 14883 3123 14909
rect 3149 14883 3175 14909
rect 20889 14883 20915 14909
rect 20941 14883 20967 14909
rect 20993 14883 21019 14909
rect 21045 14883 21071 14909
rect 21097 14883 21123 14909
rect 21149 14883 21175 14909
rect 1029 14491 1055 14517
rect 1081 14491 1107 14517
rect 1133 14491 1159 14517
rect 1185 14491 1211 14517
rect 1237 14491 1263 14517
rect 1289 14491 1315 14517
rect 19029 14491 19055 14517
rect 19081 14491 19107 14517
rect 19133 14491 19159 14517
rect 19185 14491 19211 14517
rect 19237 14491 19263 14517
rect 19289 14491 19315 14517
rect 2889 14099 2915 14125
rect 2941 14099 2967 14125
rect 2993 14099 3019 14125
rect 3045 14099 3071 14125
rect 3097 14099 3123 14125
rect 3149 14099 3175 14125
rect 20889 14099 20915 14125
rect 20941 14099 20967 14125
rect 20993 14099 21019 14125
rect 21045 14099 21071 14125
rect 21097 14099 21123 14125
rect 21149 14099 21175 14125
rect 1029 13707 1055 13733
rect 1081 13707 1107 13733
rect 1133 13707 1159 13733
rect 1185 13707 1211 13733
rect 1237 13707 1263 13733
rect 1289 13707 1315 13733
rect 19029 13707 19055 13733
rect 19081 13707 19107 13733
rect 19133 13707 19159 13733
rect 19185 13707 19211 13733
rect 19237 13707 19263 13733
rect 19289 13707 19315 13733
rect 2889 13315 2915 13341
rect 2941 13315 2967 13341
rect 2993 13315 3019 13341
rect 3045 13315 3071 13341
rect 3097 13315 3123 13341
rect 3149 13315 3175 13341
rect 20889 13315 20915 13341
rect 20941 13315 20967 13341
rect 20993 13315 21019 13341
rect 21045 13315 21071 13341
rect 21097 13315 21123 13341
rect 21149 13315 21175 13341
rect 1029 12923 1055 12949
rect 1081 12923 1107 12949
rect 1133 12923 1159 12949
rect 1185 12923 1211 12949
rect 1237 12923 1263 12949
rect 1289 12923 1315 12949
rect 19029 12923 19055 12949
rect 19081 12923 19107 12949
rect 19133 12923 19159 12949
rect 19185 12923 19211 12949
rect 19237 12923 19263 12949
rect 19289 12923 19315 12949
rect 911 12615 937 12641
rect 2889 12531 2915 12557
rect 2941 12531 2967 12557
rect 2993 12531 3019 12557
rect 3045 12531 3071 12557
rect 3097 12531 3123 12557
rect 3149 12531 3175 12557
rect 20889 12531 20915 12557
rect 20941 12531 20967 12557
rect 20993 12531 21019 12557
rect 21045 12531 21071 12557
rect 21097 12531 21123 12557
rect 21149 12531 21175 12557
rect 1029 12139 1055 12165
rect 1081 12139 1107 12165
rect 1133 12139 1159 12165
rect 1185 12139 1211 12165
rect 1237 12139 1263 12165
rect 1289 12139 1315 12165
rect 19029 12139 19055 12165
rect 19081 12139 19107 12165
rect 19133 12139 19159 12165
rect 19185 12139 19211 12165
rect 19237 12139 19263 12165
rect 19289 12139 19315 12165
rect 2889 11747 2915 11773
rect 2941 11747 2967 11773
rect 2993 11747 3019 11773
rect 3045 11747 3071 11773
rect 3097 11747 3123 11773
rect 3149 11747 3175 11773
rect 20889 11747 20915 11773
rect 20941 11747 20967 11773
rect 20993 11747 21019 11773
rect 21045 11747 21071 11773
rect 21097 11747 21123 11773
rect 21149 11747 21175 11773
rect 1029 11355 1055 11381
rect 1081 11355 1107 11381
rect 1133 11355 1159 11381
rect 1185 11355 1211 11381
rect 1237 11355 1263 11381
rect 1289 11355 1315 11381
rect 19029 11355 19055 11381
rect 19081 11355 19107 11381
rect 19133 11355 19159 11381
rect 19185 11355 19211 11381
rect 19237 11355 19263 11381
rect 19289 11355 19315 11381
rect 2889 10963 2915 10989
rect 2941 10963 2967 10989
rect 2993 10963 3019 10989
rect 3045 10963 3071 10989
rect 3097 10963 3123 10989
rect 3149 10963 3175 10989
rect 20889 10963 20915 10989
rect 20941 10963 20967 10989
rect 20993 10963 21019 10989
rect 21045 10963 21071 10989
rect 21097 10963 21123 10989
rect 21149 10963 21175 10989
rect 1029 10571 1055 10597
rect 1081 10571 1107 10597
rect 1133 10571 1159 10597
rect 1185 10571 1211 10597
rect 1237 10571 1263 10597
rect 1289 10571 1315 10597
rect 19029 10571 19055 10597
rect 19081 10571 19107 10597
rect 19133 10571 19159 10597
rect 19185 10571 19211 10597
rect 19237 10571 19263 10597
rect 19289 10571 19315 10597
rect 2889 10179 2915 10205
rect 2941 10179 2967 10205
rect 2993 10179 3019 10205
rect 3045 10179 3071 10205
rect 3097 10179 3123 10205
rect 3149 10179 3175 10205
rect 20889 10179 20915 10205
rect 20941 10179 20967 10205
rect 20993 10179 21019 10205
rect 21045 10179 21071 10205
rect 21097 10179 21123 10205
rect 21149 10179 21175 10205
rect 1029 9787 1055 9813
rect 1081 9787 1107 9813
rect 1133 9787 1159 9813
rect 1185 9787 1211 9813
rect 1237 9787 1263 9813
rect 1289 9787 1315 9813
rect 19029 9787 19055 9813
rect 19081 9787 19107 9813
rect 19133 9787 19159 9813
rect 19185 9787 19211 9813
rect 19237 9787 19263 9813
rect 19289 9787 19315 9813
rect 2889 9395 2915 9421
rect 2941 9395 2967 9421
rect 2993 9395 3019 9421
rect 3045 9395 3071 9421
rect 3097 9395 3123 9421
rect 3149 9395 3175 9421
rect 20889 9395 20915 9421
rect 20941 9395 20967 9421
rect 20993 9395 21019 9421
rect 21045 9395 21071 9421
rect 21097 9395 21123 9421
rect 21149 9395 21175 9421
rect 1029 9003 1055 9029
rect 1081 9003 1107 9029
rect 1133 9003 1159 9029
rect 1185 9003 1211 9029
rect 1237 9003 1263 9029
rect 1289 9003 1315 9029
rect 19029 9003 19055 9029
rect 19081 9003 19107 9029
rect 19133 9003 19159 9029
rect 19185 9003 19211 9029
rect 19237 9003 19263 9029
rect 19289 9003 19315 9029
rect 2889 8611 2915 8637
rect 2941 8611 2967 8637
rect 2993 8611 3019 8637
rect 3045 8611 3071 8637
rect 3097 8611 3123 8637
rect 3149 8611 3175 8637
rect 20889 8611 20915 8637
rect 20941 8611 20967 8637
rect 20993 8611 21019 8637
rect 21045 8611 21071 8637
rect 21097 8611 21123 8637
rect 21149 8611 21175 8637
rect 1029 8219 1055 8245
rect 1081 8219 1107 8245
rect 1133 8219 1159 8245
rect 1185 8219 1211 8245
rect 1237 8219 1263 8245
rect 1289 8219 1315 8245
rect 19029 8219 19055 8245
rect 19081 8219 19107 8245
rect 19133 8219 19159 8245
rect 19185 8219 19211 8245
rect 19237 8219 19263 8245
rect 19289 8219 19315 8245
rect 2889 7827 2915 7853
rect 2941 7827 2967 7853
rect 2993 7827 3019 7853
rect 3045 7827 3071 7853
rect 3097 7827 3123 7853
rect 3149 7827 3175 7853
rect 20889 7827 20915 7853
rect 20941 7827 20967 7853
rect 20993 7827 21019 7853
rect 21045 7827 21071 7853
rect 21097 7827 21123 7853
rect 21149 7827 21175 7853
rect 1029 7435 1055 7461
rect 1081 7435 1107 7461
rect 1133 7435 1159 7461
rect 1185 7435 1211 7461
rect 1237 7435 1263 7461
rect 1289 7435 1315 7461
rect 19029 7435 19055 7461
rect 19081 7435 19107 7461
rect 19133 7435 19159 7461
rect 19185 7435 19211 7461
rect 19237 7435 19263 7461
rect 19289 7435 19315 7461
rect 2889 7043 2915 7069
rect 2941 7043 2967 7069
rect 2993 7043 3019 7069
rect 3045 7043 3071 7069
rect 3097 7043 3123 7069
rect 3149 7043 3175 7069
rect 20889 7043 20915 7069
rect 20941 7043 20967 7069
rect 20993 7043 21019 7069
rect 21045 7043 21071 7069
rect 21097 7043 21123 7069
rect 21149 7043 21175 7069
rect 1029 6651 1055 6677
rect 1081 6651 1107 6677
rect 1133 6651 1159 6677
rect 1185 6651 1211 6677
rect 1237 6651 1263 6677
rect 1289 6651 1315 6677
rect 19029 6651 19055 6677
rect 19081 6651 19107 6677
rect 19133 6651 19159 6677
rect 19185 6651 19211 6677
rect 19237 6651 19263 6677
rect 19289 6651 19315 6677
rect 2889 6259 2915 6285
rect 2941 6259 2967 6285
rect 2993 6259 3019 6285
rect 3045 6259 3071 6285
rect 3097 6259 3123 6285
rect 3149 6259 3175 6285
rect 20889 6259 20915 6285
rect 20941 6259 20967 6285
rect 20993 6259 21019 6285
rect 21045 6259 21071 6285
rect 21097 6259 21123 6285
rect 21149 6259 21175 6285
rect 16031 6063 16057 6089
rect 16255 6063 16281 6089
rect 13511 6007 13537 6033
rect 1029 5867 1055 5893
rect 1081 5867 1107 5893
rect 1133 5867 1159 5893
rect 1185 5867 1211 5893
rect 1237 5867 1263 5893
rect 1289 5867 1315 5893
rect 19029 5867 19055 5893
rect 19081 5867 19107 5893
rect 19133 5867 19159 5893
rect 19185 5867 19211 5893
rect 19237 5867 19263 5893
rect 19289 5867 19315 5893
rect 12503 5671 12529 5697
rect 12839 5671 12865 5697
rect 12895 5615 12921 5641
rect 12335 5559 12361 5585
rect 13231 5559 13257 5585
rect 2889 5475 2915 5501
rect 2941 5475 2967 5501
rect 2993 5475 3019 5501
rect 3045 5475 3071 5501
rect 3097 5475 3123 5501
rect 3149 5475 3175 5501
rect 20889 5475 20915 5501
rect 20941 5475 20967 5501
rect 20993 5475 21019 5501
rect 21045 5475 21071 5501
rect 21097 5475 21123 5501
rect 21149 5475 21175 5501
rect 11887 5391 11913 5417
rect 11719 5335 11745 5361
rect 12839 5279 12865 5305
rect 12503 5223 12529 5249
rect 14295 5223 14321 5249
rect 1029 5083 1055 5109
rect 1081 5083 1107 5109
rect 1133 5083 1159 5109
rect 1185 5083 1211 5109
rect 1237 5083 1263 5109
rect 1289 5083 1315 5109
rect 19029 5083 19055 5109
rect 19081 5083 19107 5109
rect 19133 5083 19159 5109
rect 19185 5083 19211 5109
rect 19237 5083 19263 5109
rect 19289 5083 19315 5109
rect 13343 4943 13369 4969
rect 11887 4887 11913 4913
rect 12279 4831 12305 4857
rect 13567 4775 13593 4801
rect 2889 4691 2915 4717
rect 2941 4691 2967 4717
rect 2993 4691 3019 4717
rect 3045 4691 3071 4717
rect 3097 4691 3123 4717
rect 3149 4691 3175 4717
rect 20889 4691 20915 4717
rect 20941 4691 20967 4717
rect 20993 4691 21019 4717
rect 21045 4691 21071 4717
rect 21097 4691 21123 4717
rect 21149 4691 21175 4717
rect 911 4551 937 4577
rect 1079 4495 1105 4521
rect 1359 4495 1385 4521
rect 1029 4299 1055 4325
rect 1081 4299 1107 4325
rect 1133 4299 1159 4325
rect 1185 4299 1211 4325
rect 1237 4299 1263 4325
rect 1289 4299 1315 4325
rect 19029 4299 19055 4325
rect 19081 4299 19107 4325
rect 19133 4299 19159 4325
rect 19185 4299 19211 4325
rect 19237 4299 19263 4325
rect 19289 4299 19315 4325
rect 2889 3907 2915 3933
rect 2941 3907 2967 3933
rect 2993 3907 3019 3933
rect 3045 3907 3071 3933
rect 3097 3907 3123 3933
rect 3149 3907 3175 3933
rect 20889 3907 20915 3933
rect 20941 3907 20967 3933
rect 20993 3907 21019 3933
rect 21045 3907 21071 3933
rect 21097 3907 21123 3933
rect 21149 3907 21175 3933
rect 10879 3767 10905 3793
rect 12223 3711 12249 3737
rect 12447 3711 12473 3737
rect 1029 3515 1055 3541
rect 1081 3515 1107 3541
rect 1133 3515 1159 3541
rect 1185 3515 1211 3541
rect 1237 3515 1263 3541
rect 1289 3515 1315 3541
rect 19029 3515 19055 3541
rect 19081 3515 19107 3541
rect 19133 3515 19159 3541
rect 19185 3515 19211 3541
rect 19237 3515 19263 3541
rect 19289 3515 19315 3541
rect 2889 3123 2915 3149
rect 2941 3123 2967 3149
rect 2993 3123 3019 3149
rect 3045 3123 3071 3149
rect 3097 3123 3123 3149
rect 3149 3123 3175 3149
rect 20889 3123 20915 3149
rect 20941 3123 20967 3149
rect 20993 3123 21019 3149
rect 21045 3123 21071 3149
rect 21097 3123 21123 3149
rect 21149 3123 21175 3149
rect 1029 2731 1055 2757
rect 1081 2731 1107 2757
rect 1133 2731 1159 2757
rect 1185 2731 1211 2757
rect 1237 2731 1263 2757
rect 1289 2731 1315 2757
rect 19029 2731 19055 2757
rect 19081 2731 19107 2757
rect 19133 2731 19159 2757
rect 19185 2731 19211 2757
rect 19237 2731 19263 2757
rect 19289 2731 19315 2757
rect 2889 2339 2915 2365
rect 2941 2339 2967 2365
rect 2993 2339 3019 2365
rect 3045 2339 3071 2365
rect 3097 2339 3123 2365
rect 3149 2339 3175 2365
rect 20889 2339 20915 2365
rect 20941 2339 20967 2365
rect 20993 2339 21019 2365
rect 21045 2339 21071 2365
rect 21097 2339 21123 2365
rect 21149 2339 21175 2365
rect 1029 1947 1055 1973
rect 1081 1947 1107 1973
rect 1133 1947 1159 1973
rect 1185 1947 1211 1973
rect 1237 1947 1263 1973
rect 1289 1947 1315 1973
rect 19029 1947 19055 1973
rect 19081 1947 19107 1973
rect 19133 1947 19159 1973
rect 19185 1947 19211 1973
rect 19237 1947 19263 1973
rect 19289 1947 19315 1973
rect 18607 1695 18633 1721
rect 18999 1695 19025 1721
rect 18831 1639 18857 1665
rect 2889 1555 2915 1581
rect 2941 1555 2967 1581
rect 2993 1555 3019 1581
rect 3045 1555 3071 1581
rect 3097 1555 3123 1581
rect 3149 1555 3175 1581
rect 20889 1555 20915 1581
rect 20941 1555 20967 1581
rect 20993 1555 21019 1581
rect 21045 1555 21071 1581
rect 21097 1555 21123 1581
rect 21149 1555 21175 1581
<< metal2 >>
rect 1028 23142 1316 23147
rect 1056 23114 1080 23142
rect 1108 23114 1132 23142
rect 1160 23114 1184 23142
rect 1212 23114 1236 23142
rect 1264 23114 1288 23142
rect 1028 23109 1316 23114
rect 19028 23142 19316 23147
rect 19056 23114 19080 23142
rect 19108 23114 19132 23142
rect 19160 23114 19184 23142
rect 19212 23114 19236 23142
rect 19264 23114 19288 23142
rect 19028 23109 19316 23114
rect 2888 22750 3176 22755
rect 2916 22722 2940 22750
rect 2968 22722 2992 22750
rect 3020 22722 3044 22750
rect 3072 22722 3096 22750
rect 3124 22722 3148 22750
rect 2888 22717 3176 22722
rect 20888 22750 21176 22755
rect 20916 22722 20940 22750
rect 20968 22722 20992 22750
rect 21020 22722 21044 22750
rect 21072 22722 21096 22750
rect 21124 22722 21148 22750
rect 20888 22717 21176 22722
rect 1028 22358 1316 22363
rect 1056 22330 1080 22358
rect 1108 22330 1132 22358
rect 1160 22330 1184 22358
rect 1212 22330 1236 22358
rect 1264 22330 1288 22358
rect 1028 22325 1316 22330
rect 19028 22358 19316 22363
rect 19056 22330 19080 22358
rect 19108 22330 19132 22358
rect 19160 22330 19184 22358
rect 19212 22330 19236 22358
rect 19264 22330 19288 22358
rect 19028 22325 19316 22330
rect 2888 21966 3176 21971
rect 2916 21938 2940 21966
rect 2968 21938 2992 21966
rect 3020 21938 3044 21966
rect 3072 21938 3096 21966
rect 3124 21938 3148 21966
rect 2888 21933 3176 21938
rect 20888 21966 21176 21971
rect 20916 21938 20940 21966
rect 20968 21938 20992 21966
rect 21020 21938 21044 21966
rect 21072 21938 21096 21966
rect 21124 21938 21148 21966
rect 20888 21933 21176 21938
rect 1028 21574 1316 21579
rect 1056 21546 1080 21574
rect 1108 21546 1132 21574
rect 1160 21546 1184 21574
rect 1212 21546 1236 21574
rect 1264 21546 1288 21574
rect 1028 21541 1316 21546
rect 19028 21574 19316 21579
rect 19056 21546 19080 21574
rect 19108 21546 19132 21574
rect 19160 21546 19184 21574
rect 19212 21546 19236 21574
rect 19264 21546 19288 21574
rect 19028 21541 19316 21546
rect 2888 21182 3176 21187
rect 2916 21154 2940 21182
rect 2968 21154 2992 21182
rect 3020 21154 3044 21182
rect 3072 21154 3096 21182
rect 3124 21154 3148 21182
rect 2888 21149 3176 21154
rect 20888 21182 21176 21187
rect 20916 21154 20940 21182
rect 20968 21154 20992 21182
rect 21020 21154 21044 21182
rect 21072 21154 21096 21182
rect 21124 21154 21148 21182
rect 20888 21149 21176 21154
rect 910 21041 938 21047
rect 910 21015 911 21041
rect 937 21015 938 21041
rect 910 20818 938 21015
rect 910 20785 938 20790
rect 1028 20790 1316 20795
rect 1056 20762 1080 20790
rect 1108 20762 1132 20790
rect 1160 20762 1184 20790
rect 1212 20762 1236 20790
rect 1264 20762 1288 20790
rect 1028 20757 1316 20762
rect 19028 20790 19316 20795
rect 19056 20762 19080 20790
rect 19108 20762 19132 20790
rect 19160 20762 19184 20790
rect 19212 20762 19236 20790
rect 19264 20762 19288 20790
rect 19028 20757 19316 20762
rect 2888 20398 3176 20403
rect 2916 20370 2940 20398
rect 2968 20370 2992 20398
rect 3020 20370 3044 20398
rect 3072 20370 3096 20398
rect 3124 20370 3148 20398
rect 2888 20365 3176 20370
rect 20888 20398 21176 20403
rect 20916 20370 20940 20398
rect 20968 20370 20992 20398
rect 21020 20370 21044 20398
rect 21072 20370 21096 20398
rect 21124 20370 21148 20398
rect 20888 20365 21176 20370
rect 1028 20006 1316 20011
rect 1056 19978 1080 20006
rect 1108 19978 1132 20006
rect 1160 19978 1184 20006
rect 1212 19978 1236 20006
rect 1264 19978 1288 20006
rect 1028 19973 1316 19978
rect 19028 20006 19316 20011
rect 19056 19978 19080 20006
rect 19108 19978 19132 20006
rect 19160 19978 19184 20006
rect 19212 19978 19236 20006
rect 19264 19978 19288 20006
rect 19028 19973 19316 19978
rect 2888 19614 3176 19619
rect 2916 19586 2940 19614
rect 2968 19586 2992 19614
rect 3020 19586 3044 19614
rect 3072 19586 3096 19614
rect 3124 19586 3148 19614
rect 2888 19581 3176 19586
rect 20888 19614 21176 19619
rect 20916 19586 20940 19614
rect 20968 19586 20992 19614
rect 21020 19586 21044 19614
rect 21072 19586 21096 19614
rect 21124 19586 21148 19614
rect 20888 19581 21176 19586
rect 1028 19222 1316 19227
rect 1056 19194 1080 19222
rect 1108 19194 1132 19222
rect 1160 19194 1184 19222
rect 1212 19194 1236 19222
rect 1264 19194 1288 19222
rect 1028 19189 1316 19194
rect 19028 19222 19316 19227
rect 19056 19194 19080 19222
rect 19108 19194 19132 19222
rect 19160 19194 19184 19222
rect 19212 19194 19236 19222
rect 19264 19194 19288 19222
rect 19028 19189 19316 19194
rect 2888 18830 3176 18835
rect 2916 18802 2940 18830
rect 2968 18802 2992 18830
rect 3020 18802 3044 18830
rect 3072 18802 3096 18830
rect 3124 18802 3148 18830
rect 2888 18797 3176 18802
rect 20888 18830 21176 18835
rect 20916 18802 20940 18830
rect 20968 18802 20992 18830
rect 21020 18802 21044 18830
rect 21072 18802 21096 18830
rect 21124 18802 21148 18830
rect 20888 18797 21176 18802
rect 1028 18438 1316 18443
rect 1056 18410 1080 18438
rect 1108 18410 1132 18438
rect 1160 18410 1184 18438
rect 1212 18410 1236 18438
rect 1264 18410 1288 18438
rect 1028 18405 1316 18410
rect 19028 18438 19316 18443
rect 19056 18410 19080 18438
rect 19108 18410 19132 18438
rect 19160 18410 19184 18438
rect 19212 18410 19236 18438
rect 19264 18410 19288 18438
rect 19028 18405 19316 18410
rect 2888 18046 3176 18051
rect 2916 18018 2940 18046
rect 2968 18018 2992 18046
rect 3020 18018 3044 18046
rect 3072 18018 3096 18046
rect 3124 18018 3148 18046
rect 2888 18013 3176 18018
rect 20888 18046 21176 18051
rect 20916 18018 20940 18046
rect 20968 18018 20992 18046
rect 21020 18018 21044 18046
rect 21072 18018 21096 18046
rect 21124 18018 21148 18046
rect 20888 18013 21176 18018
rect 1028 17654 1316 17659
rect 1056 17626 1080 17654
rect 1108 17626 1132 17654
rect 1160 17626 1184 17654
rect 1212 17626 1236 17654
rect 1264 17626 1288 17654
rect 1028 17621 1316 17626
rect 19028 17654 19316 17659
rect 19056 17626 19080 17654
rect 19108 17626 19132 17654
rect 19160 17626 19184 17654
rect 19212 17626 19236 17654
rect 19264 17626 19288 17654
rect 19028 17621 19316 17626
rect 2888 17262 3176 17267
rect 2916 17234 2940 17262
rect 2968 17234 2992 17262
rect 3020 17234 3044 17262
rect 3072 17234 3096 17262
rect 3124 17234 3148 17262
rect 2888 17229 3176 17234
rect 20888 17262 21176 17267
rect 20916 17234 20940 17262
rect 20968 17234 20992 17262
rect 21020 17234 21044 17262
rect 21072 17234 21096 17262
rect 21124 17234 21148 17262
rect 20888 17229 21176 17234
rect 1028 16870 1316 16875
rect 1056 16842 1080 16870
rect 1108 16842 1132 16870
rect 1160 16842 1184 16870
rect 1212 16842 1236 16870
rect 1264 16842 1288 16870
rect 1028 16837 1316 16842
rect 19028 16870 19316 16875
rect 19056 16842 19080 16870
rect 19108 16842 19132 16870
rect 19160 16842 19184 16870
rect 19212 16842 19236 16870
rect 19264 16842 19288 16870
rect 19028 16837 19316 16842
rect 2888 16478 3176 16483
rect 2916 16450 2940 16478
rect 2968 16450 2992 16478
rect 3020 16450 3044 16478
rect 3072 16450 3096 16478
rect 3124 16450 3148 16478
rect 2888 16445 3176 16450
rect 20888 16478 21176 16483
rect 20916 16450 20940 16478
rect 20968 16450 20992 16478
rect 21020 16450 21044 16478
rect 21072 16450 21096 16478
rect 21124 16450 21148 16478
rect 20888 16445 21176 16450
rect 1028 16086 1316 16091
rect 1056 16058 1080 16086
rect 1108 16058 1132 16086
rect 1160 16058 1184 16086
rect 1212 16058 1236 16086
rect 1264 16058 1288 16086
rect 1028 16053 1316 16058
rect 19028 16086 19316 16091
rect 19056 16058 19080 16086
rect 19108 16058 19132 16086
rect 19160 16058 19184 16086
rect 19212 16058 19236 16086
rect 19264 16058 19288 16086
rect 19028 16053 19316 16058
rect 2888 15694 3176 15699
rect 2916 15666 2940 15694
rect 2968 15666 2992 15694
rect 3020 15666 3044 15694
rect 3072 15666 3096 15694
rect 3124 15666 3148 15694
rect 2888 15661 3176 15666
rect 20888 15694 21176 15699
rect 20916 15666 20940 15694
rect 20968 15666 20992 15694
rect 21020 15666 21044 15694
rect 21072 15666 21096 15694
rect 21124 15666 21148 15694
rect 20888 15661 21176 15666
rect 1028 15302 1316 15307
rect 1056 15274 1080 15302
rect 1108 15274 1132 15302
rect 1160 15274 1184 15302
rect 1212 15274 1236 15302
rect 1264 15274 1288 15302
rect 1028 15269 1316 15274
rect 19028 15302 19316 15307
rect 19056 15274 19080 15302
rect 19108 15274 19132 15302
rect 19160 15274 19184 15302
rect 19212 15274 19236 15302
rect 19264 15274 19288 15302
rect 19028 15269 19316 15274
rect 2888 14910 3176 14915
rect 2916 14882 2940 14910
rect 2968 14882 2992 14910
rect 3020 14882 3044 14910
rect 3072 14882 3096 14910
rect 3124 14882 3148 14910
rect 2888 14877 3176 14882
rect 20888 14910 21176 14915
rect 20916 14882 20940 14910
rect 20968 14882 20992 14910
rect 21020 14882 21044 14910
rect 21072 14882 21096 14910
rect 21124 14882 21148 14910
rect 20888 14877 21176 14882
rect 1028 14518 1316 14523
rect 1056 14490 1080 14518
rect 1108 14490 1132 14518
rect 1160 14490 1184 14518
rect 1212 14490 1236 14518
rect 1264 14490 1288 14518
rect 1028 14485 1316 14490
rect 19028 14518 19316 14523
rect 19056 14490 19080 14518
rect 19108 14490 19132 14518
rect 19160 14490 19184 14518
rect 19212 14490 19236 14518
rect 19264 14490 19288 14518
rect 19028 14485 19316 14490
rect 2888 14126 3176 14131
rect 2916 14098 2940 14126
rect 2968 14098 2992 14126
rect 3020 14098 3044 14126
rect 3072 14098 3096 14126
rect 3124 14098 3148 14126
rect 2888 14093 3176 14098
rect 20888 14126 21176 14131
rect 20916 14098 20940 14126
rect 20968 14098 20992 14126
rect 21020 14098 21044 14126
rect 21072 14098 21096 14126
rect 21124 14098 21148 14126
rect 20888 14093 21176 14098
rect 1028 13734 1316 13739
rect 1056 13706 1080 13734
rect 1108 13706 1132 13734
rect 1160 13706 1184 13734
rect 1212 13706 1236 13734
rect 1264 13706 1288 13734
rect 1028 13701 1316 13706
rect 19028 13734 19316 13739
rect 19056 13706 19080 13734
rect 19108 13706 19132 13734
rect 19160 13706 19184 13734
rect 19212 13706 19236 13734
rect 19264 13706 19288 13734
rect 19028 13701 19316 13706
rect 2888 13342 3176 13347
rect 2916 13314 2940 13342
rect 2968 13314 2992 13342
rect 3020 13314 3044 13342
rect 3072 13314 3096 13342
rect 3124 13314 3148 13342
rect 2888 13309 3176 13314
rect 20888 13342 21176 13347
rect 20916 13314 20940 13342
rect 20968 13314 20992 13342
rect 21020 13314 21044 13342
rect 21072 13314 21096 13342
rect 21124 13314 21148 13342
rect 20888 13309 21176 13314
rect 1028 12950 1316 12955
rect 1056 12922 1080 12950
rect 1108 12922 1132 12950
rect 1160 12922 1184 12950
rect 1212 12922 1236 12950
rect 1264 12922 1288 12950
rect 1028 12917 1316 12922
rect 19028 12950 19316 12955
rect 19056 12922 19080 12950
rect 19108 12922 19132 12950
rect 19160 12922 19184 12950
rect 19212 12922 19236 12950
rect 19264 12922 19288 12950
rect 19028 12917 19316 12922
rect 910 12641 938 12647
rect 910 12615 911 12641
rect 937 12615 938 12641
rect 910 12530 938 12615
rect 2888 12558 3176 12563
rect 2916 12530 2940 12558
rect 2968 12530 2992 12558
rect 3020 12530 3044 12558
rect 3072 12530 3096 12558
rect 3124 12530 3148 12558
rect 2888 12525 3176 12530
rect 20888 12558 21176 12563
rect 20916 12530 20940 12558
rect 20968 12530 20992 12558
rect 21020 12530 21044 12558
rect 21072 12530 21096 12558
rect 21124 12530 21148 12558
rect 20888 12525 21176 12530
rect 910 12497 938 12502
rect 22246 12474 22274 12479
rect 1028 12166 1316 12171
rect 1056 12138 1080 12166
rect 1108 12138 1132 12166
rect 1160 12138 1184 12166
rect 1212 12138 1236 12166
rect 1264 12138 1288 12166
rect 1028 12133 1316 12138
rect 19028 12166 19316 12171
rect 19056 12138 19080 12166
rect 19108 12138 19132 12166
rect 19160 12138 19184 12166
rect 19212 12138 19236 12166
rect 19264 12138 19288 12166
rect 19028 12133 19316 12138
rect 2888 11774 3176 11779
rect 2916 11746 2940 11774
rect 2968 11746 2992 11774
rect 3020 11746 3044 11774
rect 3072 11746 3096 11774
rect 3124 11746 3148 11774
rect 2888 11741 3176 11746
rect 20888 11774 21176 11779
rect 20916 11746 20940 11774
rect 20968 11746 20992 11774
rect 21020 11746 21044 11774
rect 21072 11746 21096 11774
rect 21124 11746 21148 11774
rect 20888 11741 21176 11746
rect 1028 11382 1316 11387
rect 1056 11354 1080 11382
rect 1108 11354 1132 11382
rect 1160 11354 1184 11382
rect 1212 11354 1236 11382
rect 1264 11354 1288 11382
rect 1028 11349 1316 11354
rect 19028 11382 19316 11387
rect 19056 11354 19080 11382
rect 19108 11354 19132 11382
rect 19160 11354 19184 11382
rect 19212 11354 19236 11382
rect 19264 11354 19288 11382
rect 19028 11349 19316 11354
rect 2888 10990 3176 10995
rect 2916 10962 2940 10990
rect 2968 10962 2992 10990
rect 3020 10962 3044 10990
rect 3072 10962 3096 10990
rect 3124 10962 3148 10990
rect 2888 10957 3176 10962
rect 20888 10990 21176 10995
rect 20916 10962 20940 10990
rect 20968 10962 20992 10990
rect 21020 10962 21044 10990
rect 21072 10962 21096 10990
rect 21124 10962 21148 10990
rect 20888 10957 21176 10962
rect 1028 10598 1316 10603
rect 1056 10570 1080 10598
rect 1108 10570 1132 10598
rect 1160 10570 1184 10598
rect 1212 10570 1236 10598
rect 1264 10570 1288 10598
rect 1028 10565 1316 10570
rect 19028 10598 19316 10603
rect 19056 10570 19080 10598
rect 19108 10570 19132 10598
rect 19160 10570 19184 10598
rect 19212 10570 19236 10598
rect 19264 10570 19288 10598
rect 19028 10565 19316 10570
rect 2888 10206 3176 10211
rect 2916 10178 2940 10206
rect 2968 10178 2992 10206
rect 3020 10178 3044 10206
rect 3072 10178 3096 10206
rect 3124 10178 3148 10206
rect 2888 10173 3176 10178
rect 20888 10206 21176 10211
rect 20916 10178 20940 10206
rect 20968 10178 20992 10206
rect 21020 10178 21044 10206
rect 21072 10178 21096 10206
rect 21124 10178 21148 10206
rect 20888 10173 21176 10178
rect 1028 9814 1316 9819
rect 1056 9786 1080 9814
rect 1108 9786 1132 9814
rect 1160 9786 1184 9814
rect 1212 9786 1236 9814
rect 1264 9786 1288 9814
rect 1028 9781 1316 9786
rect 19028 9814 19316 9819
rect 19056 9786 19080 9814
rect 19108 9786 19132 9814
rect 19160 9786 19184 9814
rect 19212 9786 19236 9814
rect 19264 9786 19288 9814
rect 19028 9781 19316 9786
rect 2888 9422 3176 9427
rect 2916 9394 2940 9422
rect 2968 9394 2992 9422
rect 3020 9394 3044 9422
rect 3072 9394 3096 9422
rect 3124 9394 3148 9422
rect 2888 9389 3176 9394
rect 20888 9422 21176 9427
rect 20916 9394 20940 9422
rect 20968 9394 20992 9422
rect 21020 9394 21044 9422
rect 21072 9394 21096 9422
rect 21124 9394 21148 9422
rect 20888 9389 21176 9394
rect 1028 9030 1316 9035
rect 1056 9002 1080 9030
rect 1108 9002 1132 9030
rect 1160 9002 1184 9030
rect 1212 9002 1236 9030
rect 1264 9002 1288 9030
rect 1028 8997 1316 9002
rect 19028 9030 19316 9035
rect 19056 9002 19080 9030
rect 19108 9002 19132 9030
rect 19160 9002 19184 9030
rect 19212 9002 19236 9030
rect 19264 9002 19288 9030
rect 19028 8997 19316 9002
rect 2888 8638 3176 8643
rect 2916 8610 2940 8638
rect 2968 8610 2992 8638
rect 3020 8610 3044 8638
rect 3072 8610 3096 8638
rect 3124 8610 3148 8638
rect 2888 8605 3176 8610
rect 20888 8638 21176 8643
rect 20916 8610 20940 8638
rect 20968 8610 20992 8638
rect 21020 8610 21044 8638
rect 21072 8610 21096 8638
rect 21124 8610 21148 8638
rect 20888 8605 21176 8610
rect 1028 8246 1316 8251
rect 1056 8218 1080 8246
rect 1108 8218 1132 8246
rect 1160 8218 1184 8246
rect 1212 8218 1236 8246
rect 1264 8218 1288 8246
rect 1028 8213 1316 8218
rect 19028 8246 19316 8251
rect 19056 8218 19080 8246
rect 19108 8218 19132 8246
rect 19160 8218 19184 8246
rect 19212 8218 19236 8246
rect 19264 8218 19288 8246
rect 19028 8213 19316 8218
rect 2888 7854 3176 7859
rect 2916 7826 2940 7854
rect 2968 7826 2992 7854
rect 3020 7826 3044 7854
rect 3072 7826 3096 7854
rect 3124 7826 3148 7854
rect 2888 7821 3176 7826
rect 20888 7854 21176 7859
rect 20916 7826 20940 7854
rect 20968 7826 20992 7854
rect 21020 7826 21044 7854
rect 21072 7826 21096 7854
rect 21124 7826 21148 7854
rect 20888 7821 21176 7826
rect 1028 7462 1316 7467
rect 1056 7434 1080 7462
rect 1108 7434 1132 7462
rect 1160 7434 1184 7462
rect 1212 7434 1236 7462
rect 1264 7434 1288 7462
rect 1028 7429 1316 7434
rect 19028 7462 19316 7467
rect 19056 7434 19080 7462
rect 19108 7434 19132 7462
rect 19160 7434 19184 7462
rect 19212 7434 19236 7462
rect 19264 7434 19288 7462
rect 19028 7429 19316 7434
rect 2888 7070 3176 7075
rect 2916 7042 2940 7070
rect 2968 7042 2992 7070
rect 3020 7042 3044 7070
rect 3072 7042 3096 7070
rect 3124 7042 3148 7070
rect 2888 7037 3176 7042
rect 20888 7070 21176 7075
rect 20916 7042 20940 7070
rect 20968 7042 20992 7070
rect 21020 7042 21044 7070
rect 21072 7042 21096 7070
rect 21124 7042 21148 7070
rect 20888 7037 21176 7042
rect 1028 6678 1316 6683
rect 1056 6650 1080 6678
rect 1108 6650 1132 6678
rect 1160 6650 1184 6678
rect 1212 6650 1236 6678
rect 1264 6650 1288 6678
rect 1028 6645 1316 6650
rect 19028 6678 19316 6683
rect 19056 6650 19080 6678
rect 19108 6650 19132 6678
rect 19160 6650 19184 6678
rect 19212 6650 19236 6678
rect 19264 6650 19288 6678
rect 19028 6645 19316 6650
rect 2888 6286 3176 6291
rect 2916 6258 2940 6286
rect 2968 6258 2992 6286
rect 3020 6258 3044 6286
rect 3072 6258 3096 6286
rect 3124 6258 3148 6286
rect 2888 6253 3176 6258
rect 20888 6286 21176 6291
rect 20916 6258 20940 6286
rect 20968 6258 20992 6286
rect 21020 6258 21044 6286
rect 21072 6258 21096 6286
rect 21124 6258 21148 6286
rect 20888 6253 21176 6258
rect 14294 6090 14322 6095
rect 12894 6034 12922 6039
rect 1028 5894 1316 5899
rect 1056 5866 1080 5894
rect 1108 5866 1132 5894
rect 1160 5866 1184 5894
rect 1212 5866 1236 5894
rect 1264 5866 1288 5894
rect 1028 5861 1316 5866
rect 12502 5697 12530 5703
rect 12502 5671 12503 5697
rect 12529 5671 12530 5697
rect 12334 5586 12362 5591
rect 11886 5585 12362 5586
rect 11886 5559 12335 5585
rect 12361 5559 12362 5585
rect 11886 5558 12362 5559
rect 2888 5502 3176 5507
rect 2916 5474 2940 5502
rect 2968 5474 2992 5502
rect 3020 5474 3044 5502
rect 3072 5474 3096 5502
rect 3124 5474 3148 5502
rect 2888 5469 3176 5474
rect 11886 5417 11914 5558
rect 12334 5553 12362 5558
rect 12502 5586 12530 5671
rect 12502 5553 12530 5558
rect 12838 5697 12866 5703
rect 12838 5671 12839 5697
rect 12865 5671 12866 5697
rect 11886 5391 11887 5417
rect 11913 5391 11914 5417
rect 11886 5385 11914 5391
rect 12838 5418 12866 5671
rect 12894 5641 12922 6006
rect 13510 6034 13538 6039
rect 13510 5987 13538 6006
rect 12894 5615 12895 5641
rect 12921 5615 12922 5641
rect 12894 5609 12922 5615
rect 13230 5586 13258 5591
rect 13230 5539 13258 5558
rect 12838 5390 12922 5418
rect 11718 5361 11746 5367
rect 11718 5335 11719 5361
rect 11745 5335 11746 5361
rect 6286 5250 6314 5255
rect 1028 5110 1316 5115
rect 1056 5082 1080 5110
rect 1108 5082 1132 5110
rect 1160 5082 1184 5110
rect 1212 5082 1236 5110
rect 1264 5082 1288 5110
rect 1028 5077 1316 5082
rect 2888 4718 3176 4723
rect 2916 4690 2940 4718
rect 2968 4690 2992 4718
rect 3020 4690 3044 4718
rect 3072 4690 3096 4718
rect 3124 4690 3148 4718
rect 2888 4685 3176 4690
rect 910 4577 938 4583
rect 910 4551 911 4577
rect 937 4551 938 4577
rect 910 4186 938 4551
rect 1078 4522 1106 4527
rect 1078 4475 1106 4494
rect 1358 4522 1386 4527
rect 1358 4475 1386 4494
rect 1028 4326 1316 4331
rect 1056 4298 1080 4326
rect 1108 4298 1132 4326
rect 1160 4298 1184 4326
rect 1212 4298 1236 4326
rect 1264 4298 1288 4326
rect 1028 4293 1316 4298
rect 910 4153 938 4158
rect 2888 3934 3176 3939
rect 2916 3906 2940 3934
rect 2968 3906 2992 3934
rect 3020 3906 3044 3934
rect 3072 3906 3096 3934
rect 3124 3906 3148 3934
rect 2888 3901 3176 3906
rect 1028 3542 1316 3547
rect 1056 3514 1080 3542
rect 1108 3514 1132 3542
rect 1160 3514 1184 3542
rect 1212 3514 1236 3542
rect 1264 3514 1288 3542
rect 1028 3509 1316 3514
rect 2888 3150 3176 3155
rect 2916 3122 2940 3150
rect 2968 3122 2992 3150
rect 3020 3122 3044 3150
rect 3072 3122 3096 3150
rect 3124 3122 3148 3150
rect 2888 3117 3176 3122
rect 1028 2758 1316 2763
rect 1056 2730 1080 2758
rect 1108 2730 1132 2758
rect 1160 2730 1184 2758
rect 1212 2730 1236 2758
rect 1264 2730 1288 2758
rect 1028 2725 1316 2730
rect 2888 2366 3176 2371
rect 2916 2338 2940 2366
rect 2968 2338 2992 2366
rect 3020 2338 3044 2366
rect 3072 2338 3096 2366
rect 3124 2338 3148 2366
rect 2888 2333 3176 2338
rect 1028 1974 1316 1979
rect 1056 1946 1080 1974
rect 1108 1946 1132 1974
rect 1160 1946 1184 1974
rect 1212 1946 1236 1974
rect 1264 1946 1288 1974
rect 1028 1941 1316 1946
rect 2888 1582 3176 1587
rect 2916 1554 2940 1582
rect 2968 1554 2992 1582
rect 3020 1554 3044 1582
rect 3072 1554 3096 1582
rect 3124 1554 3148 1582
rect 2888 1549 3176 1554
rect 6286 240 6314 5222
rect 10878 4914 10906 4919
rect 10878 3793 10906 4886
rect 11718 4522 11746 5335
rect 12838 5305 12866 5311
rect 12838 5279 12839 5305
rect 12865 5279 12866 5305
rect 12502 5250 12530 5255
rect 12502 5203 12530 5222
rect 12838 5250 12866 5279
rect 12838 5217 12866 5222
rect 12446 5194 12474 5199
rect 11886 4914 11914 4919
rect 11886 4867 11914 4886
rect 12278 4857 12306 4863
rect 12278 4831 12279 4857
rect 12305 4831 12306 4857
rect 12278 4802 12306 4831
rect 12278 4769 12306 4774
rect 11718 4489 11746 4494
rect 10878 3767 10879 3793
rect 10905 3767 10906 3793
rect 10878 3761 10906 3767
rect 12222 3738 12250 3743
rect 12446 3738 12474 5166
rect 12894 4970 12922 5390
rect 14294 5249 14322 6062
rect 16030 6090 16058 6095
rect 16030 6043 16058 6062
rect 16254 6090 16282 6095
rect 16254 6043 16282 6062
rect 19028 5894 19316 5899
rect 19056 5866 19080 5894
rect 19108 5866 19132 5894
rect 19160 5866 19184 5894
rect 19212 5866 19236 5894
rect 19264 5866 19288 5894
rect 19028 5861 19316 5866
rect 22246 5586 22274 12446
rect 22246 5553 22274 5558
rect 20888 5502 21176 5507
rect 20916 5474 20940 5502
rect 20968 5474 20992 5502
rect 21020 5474 21044 5502
rect 21072 5474 21096 5502
rect 21124 5474 21148 5502
rect 20888 5469 21176 5474
rect 14294 5223 14295 5249
rect 14321 5223 14322 5249
rect 14294 5194 14322 5223
rect 14294 5161 14322 5166
rect 19028 5110 19316 5115
rect 19056 5082 19080 5110
rect 19108 5082 19132 5110
rect 19160 5082 19184 5110
rect 19212 5082 19236 5110
rect 19264 5082 19288 5110
rect 19028 5077 19316 5082
rect 13342 4970 13370 4975
rect 12894 4969 13370 4970
rect 12894 4943 13343 4969
rect 13369 4943 13370 4969
rect 12894 4942 13370 4943
rect 13342 4937 13370 4942
rect 13566 4802 13594 4807
rect 13566 4755 13594 4774
rect 18830 4802 18858 4807
rect 12222 3737 12474 3738
rect 12222 3711 12223 3737
rect 12249 3711 12447 3737
rect 12473 3711 12474 3737
rect 12222 3710 12474 3711
rect 12222 3705 12250 3710
rect 12446 3705 12474 3710
rect 18606 1722 18634 1727
rect 18662 1722 18690 1727
rect 18606 1721 18662 1722
rect 18606 1695 18607 1721
rect 18633 1695 18662 1721
rect 18606 1694 18662 1695
rect 18606 1689 18634 1694
rect 6188 196 6314 240
rect 18662 240 18690 1694
rect 18830 1665 18858 4774
rect 20888 4718 21176 4723
rect 20916 4690 20940 4718
rect 20968 4690 20992 4718
rect 21020 4690 21044 4718
rect 21072 4690 21096 4718
rect 21124 4690 21148 4718
rect 20888 4685 21176 4690
rect 19028 4326 19316 4331
rect 19056 4298 19080 4326
rect 19108 4298 19132 4326
rect 19160 4298 19184 4326
rect 19212 4298 19236 4326
rect 19264 4298 19288 4326
rect 19028 4293 19316 4298
rect 20888 3934 21176 3939
rect 20916 3906 20940 3934
rect 20968 3906 20992 3934
rect 21020 3906 21044 3934
rect 21072 3906 21096 3934
rect 21124 3906 21148 3934
rect 20888 3901 21176 3906
rect 19028 3542 19316 3547
rect 19056 3514 19080 3542
rect 19108 3514 19132 3542
rect 19160 3514 19184 3542
rect 19212 3514 19236 3542
rect 19264 3514 19288 3542
rect 19028 3509 19316 3514
rect 20888 3150 21176 3155
rect 20916 3122 20940 3150
rect 20968 3122 20992 3150
rect 21020 3122 21044 3150
rect 21072 3122 21096 3150
rect 21124 3122 21148 3150
rect 20888 3117 21176 3122
rect 19028 2758 19316 2763
rect 19056 2730 19080 2758
rect 19108 2730 19132 2758
rect 19160 2730 19184 2758
rect 19212 2730 19236 2758
rect 19264 2730 19288 2758
rect 19028 2725 19316 2730
rect 20888 2366 21176 2371
rect 20916 2338 20940 2366
rect 20968 2338 20992 2366
rect 21020 2338 21044 2366
rect 21072 2338 21096 2366
rect 21124 2338 21148 2366
rect 20888 2333 21176 2338
rect 19028 1974 19316 1979
rect 19056 1946 19080 1974
rect 19108 1946 19132 1974
rect 19160 1946 19184 1974
rect 19212 1946 19236 1974
rect 19264 1946 19288 1974
rect 19028 1941 19316 1946
rect 18998 1722 19026 1727
rect 18998 1675 19026 1694
rect 18830 1639 18831 1665
rect 18857 1639 18858 1665
rect 18830 1633 18858 1639
rect 20888 1582 21176 1587
rect 20916 1554 20940 1582
rect 20968 1554 20992 1582
rect 21020 1554 21044 1582
rect 21072 1554 21096 1582
rect 21124 1554 21148 1582
rect 20888 1549 21176 1554
rect 18662 196 18788 240
rect 6188 -480 6300 196
rect 18676 -480 18788 196
<< via2 >>
rect 1028 23141 1056 23142
rect 1028 23115 1029 23141
rect 1029 23115 1055 23141
rect 1055 23115 1056 23141
rect 1028 23114 1056 23115
rect 1080 23141 1108 23142
rect 1080 23115 1081 23141
rect 1081 23115 1107 23141
rect 1107 23115 1108 23141
rect 1080 23114 1108 23115
rect 1132 23141 1160 23142
rect 1132 23115 1133 23141
rect 1133 23115 1159 23141
rect 1159 23115 1160 23141
rect 1132 23114 1160 23115
rect 1184 23141 1212 23142
rect 1184 23115 1185 23141
rect 1185 23115 1211 23141
rect 1211 23115 1212 23141
rect 1184 23114 1212 23115
rect 1236 23141 1264 23142
rect 1236 23115 1237 23141
rect 1237 23115 1263 23141
rect 1263 23115 1264 23141
rect 1236 23114 1264 23115
rect 1288 23141 1316 23142
rect 1288 23115 1289 23141
rect 1289 23115 1315 23141
rect 1315 23115 1316 23141
rect 1288 23114 1316 23115
rect 19028 23141 19056 23142
rect 19028 23115 19029 23141
rect 19029 23115 19055 23141
rect 19055 23115 19056 23141
rect 19028 23114 19056 23115
rect 19080 23141 19108 23142
rect 19080 23115 19081 23141
rect 19081 23115 19107 23141
rect 19107 23115 19108 23141
rect 19080 23114 19108 23115
rect 19132 23141 19160 23142
rect 19132 23115 19133 23141
rect 19133 23115 19159 23141
rect 19159 23115 19160 23141
rect 19132 23114 19160 23115
rect 19184 23141 19212 23142
rect 19184 23115 19185 23141
rect 19185 23115 19211 23141
rect 19211 23115 19212 23141
rect 19184 23114 19212 23115
rect 19236 23141 19264 23142
rect 19236 23115 19237 23141
rect 19237 23115 19263 23141
rect 19263 23115 19264 23141
rect 19236 23114 19264 23115
rect 19288 23141 19316 23142
rect 19288 23115 19289 23141
rect 19289 23115 19315 23141
rect 19315 23115 19316 23141
rect 19288 23114 19316 23115
rect 2888 22749 2916 22750
rect 2888 22723 2889 22749
rect 2889 22723 2915 22749
rect 2915 22723 2916 22749
rect 2888 22722 2916 22723
rect 2940 22749 2968 22750
rect 2940 22723 2941 22749
rect 2941 22723 2967 22749
rect 2967 22723 2968 22749
rect 2940 22722 2968 22723
rect 2992 22749 3020 22750
rect 2992 22723 2993 22749
rect 2993 22723 3019 22749
rect 3019 22723 3020 22749
rect 2992 22722 3020 22723
rect 3044 22749 3072 22750
rect 3044 22723 3045 22749
rect 3045 22723 3071 22749
rect 3071 22723 3072 22749
rect 3044 22722 3072 22723
rect 3096 22749 3124 22750
rect 3096 22723 3097 22749
rect 3097 22723 3123 22749
rect 3123 22723 3124 22749
rect 3096 22722 3124 22723
rect 3148 22749 3176 22750
rect 3148 22723 3149 22749
rect 3149 22723 3175 22749
rect 3175 22723 3176 22749
rect 3148 22722 3176 22723
rect 20888 22749 20916 22750
rect 20888 22723 20889 22749
rect 20889 22723 20915 22749
rect 20915 22723 20916 22749
rect 20888 22722 20916 22723
rect 20940 22749 20968 22750
rect 20940 22723 20941 22749
rect 20941 22723 20967 22749
rect 20967 22723 20968 22749
rect 20940 22722 20968 22723
rect 20992 22749 21020 22750
rect 20992 22723 20993 22749
rect 20993 22723 21019 22749
rect 21019 22723 21020 22749
rect 20992 22722 21020 22723
rect 21044 22749 21072 22750
rect 21044 22723 21045 22749
rect 21045 22723 21071 22749
rect 21071 22723 21072 22749
rect 21044 22722 21072 22723
rect 21096 22749 21124 22750
rect 21096 22723 21097 22749
rect 21097 22723 21123 22749
rect 21123 22723 21124 22749
rect 21096 22722 21124 22723
rect 21148 22749 21176 22750
rect 21148 22723 21149 22749
rect 21149 22723 21175 22749
rect 21175 22723 21176 22749
rect 21148 22722 21176 22723
rect 1028 22357 1056 22358
rect 1028 22331 1029 22357
rect 1029 22331 1055 22357
rect 1055 22331 1056 22357
rect 1028 22330 1056 22331
rect 1080 22357 1108 22358
rect 1080 22331 1081 22357
rect 1081 22331 1107 22357
rect 1107 22331 1108 22357
rect 1080 22330 1108 22331
rect 1132 22357 1160 22358
rect 1132 22331 1133 22357
rect 1133 22331 1159 22357
rect 1159 22331 1160 22357
rect 1132 22330 1160 22331
rect 1184 22357 1212 22358
rect 1184 22331 1185 22357
rect 1185 22331 1211 22357
rect 1211 22331 1212 22357
rect 1184 22330 1212 22331
rect 1236 22357 1264 22358
rect 1236 22331 1237 22357
rect 1237 22331 1263 22357
rect 1263 22331 1264 22357
rect 1236 22330 1264 22331
rect 1288 22357 1316 22358
rect 1288 22331 1289 22357
rect 1289 22331 1315 22357
rect 1315 22331 1316 22357
rect 1288 22330 1316 22331
rect 19028 22357 19056 22358
rect 19028 22331 19029 22357
rect 19029 22331 19055 22357
rect 19055 22331 19056 22357
rect 19028 22330 19056 22331
rect 19080 22357 19108 22358
rect 19080 22331 19081 22357
rect 19081 22331 19107 22357
rect 19107 22331 19108 22357
rect 19080 22330 19108 22331
rect 19132 22357 19160 22358
rect 19132 22331 19133 22357
rect 19133 22331 19159 22357
rect 19159 22331 19160 22357
rect 19132 22330 19160 22331
rect 19184 22357 19212 22358
rect 19184 22331 19185 22357
rect 19185 22331 19211 22357
rect 19211 22331 19212 22357
rect 19184 22330 19212 22331
rect 19236 22357 19264 22358
rect 19236 22331 19237 22357
rect 19237 22331 19263 22357
rect 19263 22331 19264 22357
rect 19236 22330 19264 22331
rect 19288 22357 19316 22358
rect 19288 22331 19289 22357
rect 19289 22331 19315 22357
rect 19315 22331 19316 22357
rect 19288 22330 19316 22331
rect 2888 21965 2916 21966
rect 2888 21939 2889 21965
rect 2889 21939 2915 21965
rect 2915 21939 2916 21965
rect 2888 21938 2916 21939
rect 2940 21965 2968 21966
rect 2940 21939 2941 21965
rect 2941 21939 2967 21965
rect 2967 21939 2968 21965
rect 2940 21938 2968 21939
rect 2992 21965 3020 21966
rect 2992 21939 2993 21965
rect 2993 21939 3019 21965
rect 3019 21939 3020 21965
rect 2992 21938 3020 21939
rect 3044 21965 3072 21966
rect 3044 21939 3045 21965
rect 3045 21939 3071 21965
rect 3071 21939 3072 21965
rect 3044 21938 3072 21939
rect 3096 21965 3124 21966
rect 3096 21939 3097 21965
rect 3097 21939 3123 21965
rect 3123 21939 3124 21965
rect 3096 21938 3124 21939
rect 3148 21965 3176 21966
rect 3148 21939 3149 21965
rect 3149 21939 3175 21965
rect 3175 21939 3176 21965
rect 3148 21938 3176 21939
rect 20888 21965 20916 21966
rect 20888 21939 20889 21965
rect 20889 21939 20915 21965
rect 20915 21939 20916 21965
rect 20888 21938 20916 21939
rect 20940 21965 20968 21966
rect 20940 21939 20941 21965
rect 20941 21939 20967 21965
rect 20967 21939 20968 21965
rect 20940 21938 20968 21939
rect 20992 21965 21020 21966
rect 20992 21939 20993 21965
rect 20993 21939 21019 21965
rect 21019 21939 21020 21965
rect 20992 21938 21020 21939
rect 21044 21965 21072 21966
rect 21044 21939 21045 21965
rect 21045 21939 21071 21965
rect 21071 21939 21072 21965
rect 21044 21938 21072 21939
rect 21096 21965 21124 21966
rect 21096 21939 21097 21965
rect 21097 21939 21123 21965
rect 21123 21939 21124 21965
rect 21096 21938 21124 21939
rect 21148 21965 21176 21966
rect 21148 21939 21149 21965
rect 21149 21939 21175 21965
rect 21175 21939 21176 21965
rect 21148 21938 21176 21939
rect 1028 21573 1056 21574
rect 1028 21547 1029 21573
rect 1029 21547 1055 21573
rect 1055 21547 1056 21573
rect 1028 21546 1056 21547
rect 1080 21573 1108 21574
rect 1080 21547 1081 21573
rect 1081 21547 1107 21573
rect 1107 21547 1108 21573
rect 1080 21546 1108 21547
rect 1132 21573 1160 21574
rect 1132 21547 1133 21573
rect 1133 21547 1159 21573
rect 1159 21547 1160 21573
rect 1132 21546 1160 21547
rect 1184 21573 1212 21574
rect 1184 21547 1185 21573
rect 1185 21547 1211 21573
rect 1211 21547 1212 21573
rect 1184 21546 1212 21547
rect 1236 21573 1264 21574
rect 1236 21547 1237 21573
rect 1237 21547 1263 21573
rect 1263 21547 1264 21573
rect 1236 21546 1264 21547
rect 1288 21573 1316 21574
rect 1288 21547 1289 21573
rect 1289 21547 1315 21573
rect 1315 21547 1316 21573
rect 1288 21546 1316 21547
rect 19028 21573 19056 21574
rect 19028 21547 19029 21573
rect 19029 21547 19055 21573
rect 19055 21547 19056 21573
rect 19028 21546 19056 21547
rect 19080 21573 19108 21574
rect 19080 21547 19081 21573
rect 19081 21547 19107 21573
rect 19107 21547 19108 21573
rect 19080 21546 19108 21547
rect 19132 21573 19160 21574
rect 19132 21547 19133 21573
rect 19133 21547 19159 21573
rect 19159 21547 19160 21573
rect 19132 21546 19160 21547
rect 19184 21573 19212 21574
rect 19184 21547 19185 21573
rect 19185 21547 19211 21573
rect 19211 21547 19212 21573
rect 19184 21546 19212 21547
rect 19236 21573 19264 21574
rect 19236 21547 19237 21573
rect 19237 21547 19263 21573
rect 19263 21547 19264 21573
rect 19236 21546 19264 21547
rect 19288 21573 19316 21574
rect 19288 21547 19289 21573
rect 19289 21547 19315 21573
rect 19315 21547 19316 21573
rect 19288 21546 19316 21547
rect 2888 21181 2916 21182
rect 2888 21155 2889 21181
rect 2889 21155 2915 21181
rect 2915 21155 2916 21181
rect 2888 21154 2916 21155
rect 2940 21181 2968 21182
rect 2940 21155 2941 21181
rect 2941 21155 2967 21181
rect 2967 21155 2968 21181
rect 2940 21154 2968 21155
rect 2992 21181 3020 21182
rect 2992 21155 2993 21181
rect 2993 21155 3019 21181
rect 3019 21155 3020 21181
rect 2992 21154 3020 21155
rect 3044 21181 3072 21182
rect 3044 21155 3045 21181
rect 3045 21155 3071 21181
rect 3071 21155 3072 21181
rect 3044 21154 3072 21155
rect 3096 21181 3124 21182
rect 3096 21155 3097 21181
rect 3097 21155 3123 21181
rect 3123 21155 3124 21181
rect 3096 21154 3124 21155
rect 3148 21181 3176 21182
rect 3148 21155 3149 21181
rect 3149 21155 3175 21181
rect 3175 21155 3176 21181
rect 3148 21154 3176 21155
rect 20888 21181 20916 21182
rect 20888 21155 20889 21181
rect 20889 21155 20915 21181
rect 20915 21155 20916 21181
rect 20888 21154 20916 21155
rect 20940 21181 20968 21182
rect 20940 21155 20941 21181
rect 20941 21155 20967 21181
rect 20967 21155 20968 21181
rect 20940 21154 20968 21155
rect 20992 21181 21020 21182
rect 20992 21155 20993 21181
rect 20993 21155 21019 21181
rect 21019 21155 21020 21181
rect 20992 21154 21020 21155
rect 21044 21181 21072 21182
rect 21044 21155 21045 21181
rect 21045 21155 21071 21181
rect 21071 21155 21072 21181
rect 21044 21154 21072 21155
rect 21096 21181 21124 21182
rect 21096 21155 21097 21181
rect 21097 21155 21123 21181
rect 21123 21155 21124 21181
rect 21096 21154 21124 21155
rect 21148 21181 21176 21182
rect 21148 21155 21149 21181
rect 21149 21155 21175 21181
rect 21175 21155 21176 21181
rect 21148 21154 21176 21155
rect 910 20790 938 20818
rect 1028 20789 1056 20790
rect 1028 20763 1029 20789
rect 1029 20763 1055 20789
rect 1055 20763 1056 20789
rect 1028 20762 1056 20763
rect 1080 20789 1108 20790
rect 1080 20763 1081 20789
rect 1081 20763 1107 20789
rect 1107 20763 1108 20789
rect 1080 20762 1108 20763
rect 1132 20789 1160 20790
rect 1132 20763 1133 20789
rect 1133 20763 1159 20789
rect 1159 20763 1160 20789
rect 1132 20762 1160 20763
rect 1184 20789 1212 20790
rect 1184 20763 1185 20789
rect 1185 20763 1211 20789
rect 1211 20763 1212 20789
rect 1184 20762 1212 20763
rect 1236 20789 1264 20790
rect 1236 20763 1237 20789
rect 1237 20763 1263 20789
rect 1263 20763 1264 20789
rect 1236 20762 1264 20763
rect 1288 20789 1316 20790
rect 1288 20763 1289 20789
rect 1289 20763 1315 20789
rect 1315 20763 1316 20789
rect 1288 20762 1316 20763
rect 19028 20789 19056 20790
rect 19028 20763 19029 20789
rect 19029 20763 19055 20789
rect 19055 20763 19056 20789
rect 19028 20762 19056 20763
rect 19080 20789 19108 20790
rect 19080 20763 19081 20789
rect 19081 20763 19107 20789
rect 19107 20763 19108 20789
rect 19080 20762 19108 20763
rect 19132 20789 19160 20790
rect 19132 20763 19133 20789
rect 19133 20763 19159 20789
rect 19159 20763 19160 20789
rect 19132 20762 19160 20763
rect 19184 20789 19212 20790
rect 19184 20763 19185 20789
rect 19185 20763 19211 20789
rect 19211 20763 19212 20789
rect 19184 20762 19212 20763
rect 19236 20789 19264 20790
rect 19236 20763 19237 20789
rect 19237 20763 19263 20789
rect 19263 20763 19264 20789
rect 19236 20762 19264 20763
rect 19288 20789 19316 20790
rect 19288 20763 19289 20789
rect 19289 20763 19315 20789
rect 19315 20763 19316 20789
rect 19288 20762 19316 20763
rect 2888 20397 2916 20398
rect 2888 20371 2889 20397
rect 2889 20371 2915 20397
rect 2915 20371 2916 20397
rect 2888 20370 2916 20371
rect 2940 20397 2968 20398
rect 2940 20371 2941 20397
rect 2941 20371 2967 20397
rect 2967 20371 2968 20397
rect 2940 20370 2968 20371
rect 2992 20397 3020 20398
rect 2992 20371 2993 20397
rect 2993 20371 3019 20397
rect 3019 20371 3020 20397
rect 2992 20370 3020 20371
rect 3044 20397 3072 20398
rect 3044 20371 3045 20397
rect 3045 20371 3071 20397
rect 3071 20371 3072 20397
rect 3044 20370 3072 20371
rect 3096 20397 3124 20398
rect 3096 20371 3097 20397
rect 3097 20371 3123 20397
rect 3123 20371 3124 20397
rect 3096 20370 3124 20371
rect 3148 20397 3176 20398
rect 3148 20371 3149 20397
rect 3149 20371 3175 20397
rect 3175 20371 3176 20397
rect 3148 20370 3176 20371
rect 20888 20397 20916 20398
rect 20888 20371 20889 20397
rect 20889 20371 20915 20397
rect 20915 20371 20916 20397
rect 20888 20370 20916 20371
rect 20940 20397 20968 20398
rect 20940 20371 20941 20397
rect 20941 20371 20967 20397
rect 20967 20371 20968 20397
rect 20940 20370 20968 20371
rect 20992 20397 21020 20398
rect 20992 20371 20993 20397
rect 20993 20371 21019 20397
rect 21019 20371 21020 20397
rect 20992 20370 21020 20371
rect 21044 20397 21072 20398
rect 21044 20371 21045 20397
rect 21045 20371 21071 20397
rect 21071 20371 21072 20397
rect 21044 20370 21072 20371
rect 21096 20397 21124 20398
rect 21096 20371 21097 20397
rect 21097 20371 21123 20397
rect 21123 20371 21124 20397
rect 21096 20370 21124 20371
rect 21148 20397 21176 20398
rect 21148 20371 21149 20397
rect 21149 20371 21175 20397
rect 21175 20371 21176 20397
rect 21148 20370 21176 20371
rect 1028 20005 1056 20006
rect 1028 19979 1029 20005
rect 1029 19979 1055 20005
rect 1055 19979 1056 20005
rect 1028 19978 1056 19979
rect 1080 20005 1108 20006
rect 1080 19979 1081 20005
rect 1081 19979 1107 20005
rect 1107 19979 1108 20005
rect 1080 19978 1108 19979
rect 1132 20005 1160 20006
rect 1132 19979 1133 20005
rect 1133 19979 1159 20005
rect 1159 19979 1160 20005
rect 1132 19978 1160 19979
rect 1184 20005 1212 20006
rect 1184 19979 1185 20005
rect 1185 19979 1211 20005
rect 1211 19979 1212 20005
rect 1184 19978 1212 19979
rect 1236 20005 1264 20006
rect 1236 19979 1237 20005
rect 1237 19979 1263 20005
rect 1263 19979 1264 20005
rect 1236 19978 1264 19979
rect 1288 20005 1316 20006
rect 1288 19979 1289 20005
rect 1289 19979 1315 20005
rect 1315 19979 1316 20005
rect 1288 19978 1316 19979
rect 19028 20005 19056 20006
rect 19028 19979 19029 20005
rect 19029 19979 19055 20005
rect 19055 19979 19056 20005
rect 19028 19978 19056 19979
rect 19080 20005 19108 20006
rect 19080 19979 19081 20005
rect 19081 19979 19107 20005
rect 19107 19979 19108 20005
rect 19080 19978 19108 19979
rect 19132 20005 19160 20006
rect 19132 19979 19133 20005
rect 19133 19979 19159 20005
rect 19159 19979 19160 20005
rect 19132 19978 19160 19979
rect 19184 20005 19212 20006
rect 19184 19979 19185 20005
rect 19185 19979 19211 20005
rect 19211 19979 19212 20005
rect 19184 19978 19212 19979
rect 19236 20005 19264 20006
rect 19236 19979 19237 20005
rect 19237 19979 19263 20005
rect 19263 19979 19264 20005
rect 19236 19978 19264 19979
rect 19288 20005 19316 20006
rect 19288 19979 19289 20005
rect 19289 19979 19315 20005
rect 19315 19979 19316 20005
rect 19288 19978 19316 19979
rect 2888 19613 2916 19614
rect 2888 19587 2889 19613
rect 2889 19587 2915 19613
rect 2915 19587 2916 19613
rect 2888 19586 2916 19587
rect 2940 19613 2968 19614
rect 2940 19587 2941 19613
rect 2941 19587 2967 19613
rect 2967 19587 2968 19613
rect 2940 19586 2968 19587
rect 2992 19613 3020 19614
rect 2992 19587 2993 19613
rect 2993 19587 3019 19613
rect 3019 19587 3020 19613
rect 2992 19586 3020 19587
rect 3044 19613 3072 19614
rect 3044 19587 3045 19613
rect 3045 19587 3071 19613
rect 3071 19587 3072 19613
rect 3044 19586 3072 19587
rect 3096 19613 3124 19614
rect 3096 19587 3097 19613
rect 3097 19587 3123 19613
rect 3123 19587 3124 19613
rect 3096 19586 3124 19587
rect 3148 19613 3176 19614
rect 3148 19587 3149 19613
rect 3149 19587 3175 19613
rect 3175 19587 3176 19613
rect 3148 19586 3176 19587
rect 20888 19613 20916 19614
rect 20888 19587 20889 19613
rect 20889 19587 20915 19613
rect 20915 19587 20916 19613
rect 20888 19586 20916 19587
rect 20940 19613 20968 19614
rect 20940 19587 20941 19613
rect 20941 19587 20967 19613
rect 20967 19587 20968 19613
rect 20940 19586 20968 19587
rect 20992 19613 21020 19614
rect 20992 19587 20993 19613
rect 20993 19587 21019 19613
rect 21019 19587 21020 19613
rect 20992 19586 21020 19587
rect 21044 19613 21072 19614
rect 21044 19587 21045 19613
rect 21045 19587 21071 19613
rect 21071 19587 21072 19613
rect 21044 19586 21072 19587
rect 21096 19613 21124 19614
rect 21096 19587 21097 19613
rect 21097 19587 21123 19613
rect 21123 19587 21124 19613
rect 21096 19586 21124 19587
rect 21148 19613 21176 19614
rect 21148 19587 21149 19613
rect 21149 19587 21175 19613
rect 21175 19587 21176 19613
rect 21148 19586 21176 19587
rect 1028 19221 1056 19222
rect 1028 19195 1029 19221
rect 1029 19195 1055 19221
rect 1055 19195 1056 19221
rect 1028 19194 1056 19195
rect 1080 19221 1108 19222
rect 1080 19195 1081 19221
rect 1081 19195 1107 19221
rect 1107 19195 1108 19221
rect 1080 19194 1108 19195
rect 1132 19221 1160 19222
rect 1132 19195 1133 19221
rect 1133 19195 1159 19221
rect 1159 19195 1160 19221
rect 1132 19194 1160 19195
rect 1184 19221 1212 19222
rect 1184 19195 1185 19221
rect 1185 19195 1211 19221
rect 1211 19195 1212 19221
rect 1184 19194 1212 19195
rect 1236 19221 1264 19222
rect 1236 19195 1237 19221
rect 1237 19195 1263 19221
rect 1263 19195 1264 19221
rect 1236 19194 1264 19195
rect 1288 19221 1316 19222
rect 1288 19195 1289 19221
rect 1289 19195 1315 19221
rect 1315 19195 1316 19221
rect 1288 19194 1316 19195
rect 19028 19221 19056 19222
rect 19028 19195 19029 19221
rect 19029 19195 19055 19221
rect 19055 19195 19056 19221
rect 19028 19194 19056 19195
rect 19080 19221 19108 19222
rect 19080 19195 19081 19221
rect 19081 19195 19107 19221
rect 19107 19195 19108 19221
rect 19080 19194 19108 19195
rect 19132 19221 19160 19222
rect 19132 19195 19133 19221
rect 19133 19195 19159 19221
rect 19159 19195 19160 19221
rect 19132 19194 19160 19195
rect 19184 19221 19212 19222
rect 19184 19195 19185 19221
rect 19185 19195 19211 19221
rect 19211 19195 19212 19221
rect 19184 19194 19212 19195
rect 19236 19221 19264 19222
rect 19236 19195 19237 19221
rect 19237 19195 19263 19221
rect 19263 19195 19264 19221
rect 19236 19194 19264 19195
rect 19288 19221 19316 19222
rect 19288 19195 19289 19221
rect 19289 19195 19315 19221
rect 19315 19195 19316 19221
rect 19288 19194 19316 19195
rect 2888 18829 2916 18830
rect 2888 18803 2889 18829
rect 2889 18803 2915 18829
rect 2915 18803 2916 18829
rect 2888 18802 2916 18803
rect 2940 18829 2968 18830
rect 2940 18803 2941 18829
rect 2941 18803 2967 18829
rect 2967 18803 2968 18829
rect 2940 18802 2968 18803
rect 2992 18829 3020 18830
rect 2992 18803 2993 18829
rect 2993 18803 3019 18829
rect 3019 18803 3020 18829
rect 2992 18802 3020 18803
rect 3044 18829 3072 18830
rect 3044 18803 3045 18829
rect 3045 18803 3071 18829
rect 3071 18803 3072 18829
rect 3044 18802 3072 18803
rect 3096 18829 3124 18830
rect 3096 18803 3097 18829
rect 3097 18803 3123 18829
rect 3123 18803 3124 18829
rect 3096 18802 3124 18803
rect 3148 18829 3176 18830
rect 3148 18803 3149 18829
rect 3149 18803 3175 18829
rect 3175 18803 3176 18829
rect 3148 18802 3176 18803
rect 20888 18829 20916 18830
rect 20888 18803 20889 18829
rect 20889 18803 20915 18829
rect 20915 18803 20916 18829
rect 20888 18802 20916 18803
rect 20940 18829 20968 18830
rect 20940 18803 20941 18829
rect 20941 18803 20967 18829
rect 20967 18803 20968 18829
rect 20940 18802 20968 18803
rect 20992 18829 21020 18830
rect 20992 18803 20993 18829
rect 20993 18803 21019 18829
rect 21019 18803 21020 18829
rect 20992 18802 21020 18803
rect 21044 18829 21072 18830
rect 21044 18803 21045 18829
rect 21045 18803 21071 18829
rect 21071 18803 21072 18829
rect 21044 18802 21072 18803
rect 21096 18829 21124 18830
rect 21096 18803 21097 18829
rect 21097 18803 21123 18829
rect 21123 18803 21124 18829
rect 21096 18802 21124 18803
rect 21148 18829 21176 18830
rect 21148 18803 21149 18829
rect 21149 18803 21175 18829
rect 21175 18803 21176 18829
rect 21148 18802 21176 18803
rect 1028 18437 1056 18438
rect 1028 18411 1029 18437
rect 1029 18411 1055 18437
rect 1055 18411 1056 18437
rect 1028 18410 1056 18411
rect 1080 18437 1108 18438
rect 1080 18411 1081 18437
rect 1081 18411 1107 18437
rect 1107 18411 1108 18437
rect 1080 18410 1108 18411
rect 1132 18437 1160 18438
rect 1132 18411 1133 18437
rect 1133 18411 1159 18437
rect 1159 18411 1160 18437
rect 1132 18410 1160 18411
rect 1184 18437 1212 18438
rect 1184 18411 1185 18437
rect 1185 18411 1211 18437
rect 1211 18411 1212 18437
rect 1184 18410 1212 18411
rect 1236 18437 1264 18438
rect 1236 18411 1237 18437
rect 1237 18411 1263 18437
rect 1263 18411 1264 18437
rect 1236 18410 1264 18411
rect 1288 18437 1316 18438
rect 1288 18411 1289 18437
rect 1289 18411 1315 18437
rect 1315 18411 1316 18437
rect 1288 18410 1316 18411
rect 19028 18437 19056 18438
rect 19028 18411 19029 18437
rect 19029 18411 19055 18437
rect 19055 18411 19056 18437
rect 19028 18410 19056 18411
rect 19080 18437 19108 18438
rect 19080 18411 19081 18437
rect 19081 18411 19107 18437
rect 19107 18411 19108 18437
rect 19080 18410 19108 18411
rect 19132 18437 19160 18438
rect 19132 18411 19133 18437
rect 19133 18411 19159 18437
rect 19159 18411 19160 18437
rect 19132 18410 19160 18411
rect 19184 18437 19212 18438
rect 19184 18411 19185 18437
rect 19185 18411 19211 18437
rect 19211 18411 19212 18437
rect 19184 18410 19212 18411
rect 19236 18437 19264 18438
rect 19236 18411 19237 18437
rect 19237 18411 19263 18437
rect 19263 18411 19264 18437
rect 19236 18410 19264 18411
rect 19288 18437 19316 18438
rect 19288 18411 19289 18437
rect 19289 18411 19315 18437
rect 19315 18411 19316 18437
rect 19288 18410 19316 18411
rect 2888 18045 2916 18046
rect 2888 18019 2889 18045
rect 2889 18019 2915 18045
rect 2915 18019 2916 18045
rect 2888 18018 2916 18019
rect 2940 18045 2968 18046
rect 2940 18019 2941 18045
rect 2941 18019 2967 18045
rect 2967 18019 2968 18045
rect 2940 18018 2968 18019
rect 2992 18045 3020 18046
rect 2992 18019 2993 18045
rect 2993 18019 3019 18045
rect 3019 18019 3020 18045
rect 2992 18018 3020 18019
rect 3044 18045 3072 18046
rect 3044 18019 3045 18045
rect 3045 18019 3071 18045
rect 3071 18019 3072 18045
rect 3044 18018 3072 18019
rect 3096 18045 3124 18046
rect 3096 18019 3097 18045
rect 3097 18019 3123 18045
rect 3123 18019 3124 18045
rect 3096 18018 3124 18019
rect 3148 18045 3176 18046
rect 3148 18019 3149 18045
rect 3149 18019 3175 18045
rect 3175 18019 3176 18045
rect 3148 18018 3176 18019
rect 20888 18045 20916 18046
rect 20888 18019 20889 18045
rect 20889 18019 20915 18045
rect 20915 18019 20916 18045
rect 20888 18018 20916 18019
rect 20940 18045 20968 18046
rect 20940 18019 20941 18045
rect 20941 18019 20967 18045
rect 20967 18019 20968 18045
rect 20940 18018 20968 18019
rect 20992 18045 21020 18046
rect 20992 18019 20993 18045
rect 20993 18019 21019 18045
rect 21019 18019 21020 18045
rect 20992 18018 21020 18019
rect 21044 18045 21072 18046
rect 21044 18019 21045 18045
rect 21045 18019 21071 18045
rect 21071 18019 21072 18045
rect 21044 18018 21072 18019
rect 21096 18045 21124 18046
rect 21096 18019 21097 18045
rect 21097 18019 21123 18045
rect 21123 18019 21124 18045
rect 21096 18018 21124 18019
rect 21148 18045 21176 18046
rect 21148 18019 21149 18045
rect 21149 18019 21175 18045
rect 21175 18019 21176 18045
rect 21148 18018 21176 18019
rect 1028 17653 1056 17654
rect 1028 17627 1029 17653
rect 1029 17627 1055 17653
rect 1055 17627 1056 17653
rect 1028 17626 1056 17627
rect 1080 17653 1108 17654
rect 1080 17627 1081 17653
rect 1081 17627 1107 17653
rect 1107 17627 1108 17653
rect 1080 17626 1108 17627
rect 1132 17653 1160 17654
rect 1132 17627 1133 17653
rect 1133 17627 1159 17653
rect 1159 17627 1160 17653
rect 1132 17626 1160 17627
rect 1184 17653 1212 17654
rect 1184 17627 1185 17653
rect 1185 17627 1211 17653
rect 1211 17627 1212 17653
rect 1184 17626 1212 17627
rect 1236 17653 1264 17654
rect 1236 17627 1237 17653
rect 1237 17627 1263 17653
rect 1263 17627 1264 17653
rect 1236 17626 1264 17627
rect 1288 17653 1316 17654
rect 1288 17627 1289 17653
rect 1289 17627 1315 17653
rect 1315 17627 1316 17653
rect 1288 17626 1316 17627
rect 19028 17653 19056 17654
rect 19028 17627 19029 17653
rect 19029 17627 19055 17653
rect 19055 17627 19056 17653
rect 19028 17626 19056 17627
rect 19080 17653 19108 17654
rect 19080 17627 19081 17653
rect 19081 17627 19107 17653
rect 19107 17627 19108 17653
rect 19080 17626 19108 17627
rect 19132 17653 19160 17654
rect 19132 17627 19133 17653
rect 19133 17627 19159 17653
rect 19159 17627 19160 17653
rect 19132 17626 19160 17627
rect 19184 17653 19212 17654
rect 19184 17627 19185 17653
rect 19185 17627 19211 17653
rect 19211 17627 19212 17653
rect 19184 17626 19212 17627
rect 19236 17653 19264 17654
rect 19236 17627 19237 17653
rect 19237 17627 19263 17653
rect 19263 17627 19264 17653
rect 19236 17626 19264 17627
rect 19288 17653 19316 17654
rect 19288 17627 19289 17653
rect 19289 17627 19315 17653
rect 19315 17627 19316 17653
rect 19288 17626 19316 17627
rect 2888 17261 2916 17262
rect 2888 17235 2889 17261
rect 2889 17235 2915 17261
rect 2915 17235 2916 17261
rect 2888 17234 2916 17235
rect 2940 17261 2968 17262
rect 2940 17235 2941 17261
rect 2941 17235 2967 17261
rect 2967 17235 2968 17261
rect 2940 17234 2968 17235
rect 2992 17261 3020 17262
rect 2992 17235 2993 17261
rect 2993 17235 3019 17261
rect 3019 17235 3020 17261
rect 2992 17234 3020 17235
rect 3044 17261 3072 17262
rect 3044 17235 3045 17261
rect 3045 17235 3071 17261
rect 3071 17235 3072 17261
rect 3044 17234 3072 17235
rect 3096 17261 3124 17262
rect 3096 17235 3097 17261
rect 3097 17235 3123 17261
rect 3123 17235 3124 17261
rect 3096 17234 3124 17235
rect 3148 17261 3176 17262
rect 3148 17235 3149 17261
rect 3149 17235 3175 17261
rect 3175 17235 3176 17261
rect 3148 17234 3176 17235
rect 20888 17261 20916 17262
rect 20888 17235 20889 17261
rect 20889 17235 20915 17261
rect 20915 17235 20916 17261
rect 20888 17234 20916 17235
rect 20940 17261 20968 17262
rect 20940 17235 20941 17261
rect 20941 17235 20967 17261
rect 20967 17235 20968 17261
rect 20940 17234 20968 17235
rect 20992 17261 21020 17262
rect 20992 17235 20993 17261
rect 20993 17235 21019 17261
rect 21019 17235 21020 17261
rect 20992 17234 21020 17235
rect 21044 17261 21072 17262
rect 21044 17235 21045 17261
rect 21045 17235 21071 17261
rect 21071 17235 21072 17261
rect 21044 17234 21072 17235
rect 21096 17261 21124 17262
rect 21096 17235 21097 17261
rect 21097 17235 21123 17261
rect 21123 17235 21124 17261
rect 21096 17234 21124 17235
rect 21148 17261 21176 17262
rect 21148 17235 21149 17261
rect 21149 17235 21175 17261
rect 21175 17235 21176 17261
rect 21148 17234 21176 17235
rect 1028 16869 1056 16870
rect 1028 16843 1029 16869
rect 1029 16843 1055 16869
rect 1055 16843 1056 16869
rect 1028 16842 1056 16843
rect 1080 16869 1108 16870
rect 1080 16843 1081 16869
rect 1081 16843 1107 16869
rect 1107 16843 1108 16869
rect 1080 16842 1108 16843
rect 1132 16869 1160 16870
rect 1132 16843 1133 16869
rect 1133 16843 1159 16869
rect 1159 16843 1160 16869
rect 1132 16842 1160 16843
rect 1184 16869 1212 16870
rect 1184 16843 1185 16869
rect 1185 16843 1211 16869
rect 1211 16843 1212 16869
rect 1184 16842 1212 16843
rect 1236 16869 1264 16870
rect 1236 16843 1237 16869
rect 1237 16843 1263 16869
rect 1263 16843 1264 16869
rect 1236 16842 1264 16843
rect 1288 16869 1316 16870
rect 1288 16843 1289 16869
rect 1289 16843 1315 16869
rect 1315 16843 1316 16869
rect 1288 16842 1316 16843
rect 19028 16869 19056 16870
rect 19028 16843 19029 16869
rect 19029 16843 19055 16869
rect 19055 16843 19056 16869
rect 19028 16842 19056 16843
rect 19080 16869 19108 16870
rect 19080 16843 19081 16869
rect 19081 16843 19107 16869
rect 19107 16843 19108 16869
rect 19080 16842 19108 16843
rect 19132 16869 19160 16870
rect 19132 16843 19133 16869
rect 19133 16843 19159 16869
rect 19159 16843 19160 16869
rect 19132 16842 19160 16843
rect 19184 16869 19212 16870
rect 19184 16843 19185 16869
rect 19185 16843 19211 16869
rect 19211 16843 19212 16869
rect 19184 16842 19212 16843
rect 19236 16869 19264 16870
rect 19236 16843 19237 16869
rect 19237 16843 19263 16869
rect 19263 16843 19264 16869
rect 19236 16842 19264 16843
rect 19288 16869 19316 16870
rect 19288 16843 19289 16869
rect 19289 16843 19315 16869
rect 19315 16843 19316 16869
rect 19288 16842 19316 16843
rect 2888 16477 2916 16478
rect 2888 16451 2889 16477
rect 2889 16451 2915 16477
rect 2915 16451 2916 16477
rect 2888 16450 2916 16451
rect 2940 16477 2968 16478
rect 2940 16451 2941 16477
rect 2941 16451 2967 16477
rect 2967 16451 2968 16477
rect 2940 16450 2968 16451
rect 2992 16477 3020 16478
rect 2992 16451 2993 16477
rect 2993 16451 3019 16477
rect 3019 16451 3020 16477
rect 2992 16450 3020 16451
rect 3044 16477 3072 16478
rect 3044 16451 3045 16477
rect 3045 16451 3071 16477
rect 3071 16451 3072 16477
rect 3044 16450 3072 16451
rect 3096 16477 3124 16478
rect 3096 16451 3097 16477
rect 3097 16451 3123 16477
rect 3123 16451 3124 16477
rect 3096 16450 3124 16451
rect 3148 16477 3176 16478
rect 3148 16451 3149 16477
rect 3149 16451 3175 16477
rect 3175 16451 3176 16477
rect 3148 16450 3176 16451
rect 20888 16477 20916 16478
rect 20888 16451 20889 16477
rect 20889 16451 20915 16477
rect 20915 16451 20916 16477
rect 20888 16450 20916 16451
rect 20940 16477 20968 16478
rect 20940 16451 20941 16477
rect 20941 16451 20967 16477
rect 20967 16451 20968 16477
rect 20940 16450 20968 16451
rect 20992 16477 21020 16478
rect 20992 16451 20993 16477
rect 20993 16451 21019 16477
rect 21019 16451 21020 16477
rect 20992 16450 21020 16451
rect 21044 16477 21072 16478
rect 21044 16451 21045 16477
rect 21045 16451 21071 16477
rect 21071 16451 21072 16477
rect 21044 16450 21072 16451
rect 21096 16477 21124 16478
rect 21096 16451 21097 16477
rect 21097 16451 21123 16477
rect 21123 16451 21124 16477
rect 21096 16450 21124 16451
rect 21148 16477 21176 16478
rect 21148 16451 21149 16477
rect 21149 16451 21175 16477
rect 21175 16451 21176 16477
rect 21148 16450 21176 16451
rect 1028 16085 1056 16086
rect 1028 16059 1029 16085
rect 1029 16059 1055 16085
rect 1055 16059 1056 16085
rect 1028 16058 1056 16059
rect 1080 16085 1108 16086
rect 1080 16059 1081 16085
rect 1081 16059 1107 16085
rect 1107 16059 1108 16085
rect 1080 16058 1108 16059
rect 1132 16085 1160 16086
rect 1132 16059 1133 16085
rect 1133 16059 1159 16085
rect 1159 16059 1160 16085
rect 1132 16058 1160 16059
rect 1184 16085 1212 16086
rect 1184 16059 1185 16085
rect 1185 16059 1211 16085
rect 1211 16059 1212 16085
rect 1184 16058 1212 16059
rect 1236 16085 1264 16086
rect 1236 16059 1237 16085
rect 1237 16059 1263 16085
rect 1263 16059 1264 16085
rect 1236 16058 1264 16059
rect 1288 16085 1316 16086
rect 1288 16059 1289 16085
rect 1289 16059 1315 16085
rect 1315 16059 1316 16085
rect 1288 16058 1316 16059
rect 19028 16085 19056 16086
rect 19028 16059 19029 16085
rect 19029 16059 19055 16085
rect 19055 16059 19056 16085
rect 19028 16058 19056 16059
rect 19080 16085 19108 16086
rect 19080 16059 19081 16085
rect 19081 16059 19107 16085
rect 19107 16059 19108 16085
rect 19080 16058 19108 16059
rect 19132 16085 19160 16086
rect 19132 16059 19133 16085
rect 19133 16059 19159 16085
rect 19159 16059 19160 16085
rect 19132 16058 19160 16059
rect 19184 16085 19212 16086
rect 19184 16059 19185 16085
rect 19185 16059 19211 16085
rect 19211 16059 19212 16085
rect 19184 16058 19212 16059
rect 19236 16085 19264 16086
rect 19236 16059 19237 16085
rect 19237 16059 19263 16085
rect 19263 16059 19264 16085
rect 19236 16058 19264 16059
rect 19288 16085 19316 16086
rect 19288 16059 19289 16085
rect 19289 16059 19315 16085
rect 19315 16059 19316 16085
rect 19288 16058 19316 16059
rect 2888 15693 2916 15694
rect 2888 15667 2889 15693
rect 2889 15667 2915 15693
rect 2915 15667 2916 15693
rect 2888 15666 2916 15667
rect 2940 15693 2968 15694
rect 2940 15667 2941 15693
rect 2941 15667 2967 15693
rect 2967 15667 2968 15693
rect 2940 15666 2968 15667
rect 2992 15693 3020 15694
rect 2992 15667 2993 15693
rect 2993 15667 3019 15693
rect 3019 15667 3020 15693
rect 2992 15666 3020 15667
rect 3044 15693 3072 15694
rect 3044 15667 3045 15693
rect 3045 15667 3071 15693
rect 3071 15667 3072 15693
rect 3044 15666 3072 15667
rect 3096 15693 3124 15694
rect 3096 15667 3097 15693
rect 3097 15667 3123 15693
rect 3123 15667 3124 15693
rect 3096 15666 3124 15667
rect 3148 15693 3176 15694
rect 3148 15667 3149 15693
rect 3149 15667 3175 15693
rect 3175 15667 3176 15693
rect 3148 15666 3176 15667
rect 20888 15693 20916 15694
rect 20888 15667 20889 15693
rect 20889 15667 20915 15693
rect 20915 15667 20916 15693
rect 20888 15666 20916 15667
rect 20940 15693 20968 15694
rect 20940 15667 20941 15693
rect 20941 15667 20967 15693
rect 20967 15667 20968 15693
rect 20940 15666 20968 15667
rect 20992 15693 21020 15694
rect 20992 15667 20993 15693
rect 20993 15667 21019 15693
rect 21019 15667 21020 15693
rect 20992 15666 21020 15667
rect 21044 15693 21072 15694
rect 21044 15667 21045 15693
rect 21045 15667 21071 15693
rect 21071 15667 21072 15693
rect 21044 15666 21072 15667
rect 21096 15693 21124 15694
rect 21096 15667 21097 15693
rect 21097 15667 21123 15693
rect 21123 15667 21124 15693
rect 21096 15666 21124 15667
rect 21148 15693 21176 15694
rect 21148 15667 21149 15693
rect 21149 15667 21175 15693
rect 21175 15667 21176 15693
rect 21148 15666 21176 15667
rect 1028 15301 1056 15302
rect 1028 15275 1029 15301
rect 1029 15275 1055 15301
rect 1055 15275 1056 15301
rect 1028 15274 1056 15275
rect 1080 15301 1108 15302
rect 1080 15275 1081 15301
rect 1081 15275 1107 15301
rect 1107 15275 1108 15301
rect 1080 15274 1108 15275
rect 1132 15301 1160 15302
rect 1132 15275 1133 15301
rect 1133 15275 1159 15301
rect 1159 15275 1160 15301
rect 1132 15274 1160 15275
rect 1184 15301 1212 15302
rect 1184 15275 1185 15301
rect 1185 15275 1211 15301
rect 1211 15275 1212 15301
rect 1184 15274 1212 15275
rect 1236 15301 1264 15302
rect 1236 15275 1237 15301
rect 1237 15275 1263 15301
rect 1263 15275 1264 15301
rect 1236 15274 1264 15275
rect 1288 15301 1316 15302
rect 1288 15275 1289 15301
rect 1289 15275 1315 15301
rect 1315 15275 1316 15301
rect 1288 15274 1316 15275
rect 19028 15301 19056 15302
rect 19028 15275 19029 15301
rect 19029 15275 19055 15301
rect 19055 15275 19056 15301
rect 19028 15274 19056 15275
rect 19080 15301 19108 15302
rect 19080 15275 19081 15301
rect 19081 15275 19107 15301
rect 19107 15275 19108 15301
rect 19080 15274 19108 15275
rect 19132 15301 19160 15302
rect 19132 15275 19133 15301
rect 19133 15275 19159 15301
rect 19159 15275 19160 15301
rect 19132 15274 19160 15275
rect 19184 15301 19212 15302
rect 19184 15275 19185 15301
rect 19185 15275 19211 15301
rect 19211 15275 19212 15301
rect 19184 15274 19212 15275
rect 19236 15301 19264 15302
rect 19236 15275 19237 15301
rect 19237 15275 19263 15301
rect 19263 15275 19264 15301
rect 19236 15274 19264 15275
rect 19288 15301 19316 15302
rect 19288 15275 19289 15301
rect 19289 15275 19315 15301
rect 19315 15275 19316 15301
rect 19288 15274 19316 15275
rect 2888 14909 2916 14910
rect 2888 14883 2889 14909
rect 2889 14883 2915 14909
rect 2915 14883 2916 14909
rect 2888 14882 2916 14883
rect 2940 14909 2968 14910
rect 2940 14883 2941 14909
rect 2941 14883 2967 14909
rect 2967 14883 2968 14909
rect 2940 14882 2968 14883
rect 2992 14909 3020 14910
rect 2992 14883 2993 14909
rect 2993 14883 3019 14909
rect 3019 14883 3020 14909
rect 2992 14882 3020 14883
rect 3044 14909 3072 14910
rect 3044 14883 3045 14909
rect 3045 14883 3071 14909
rect 3071 14883 3072 14909
rect 3044 14882 3072 14883
rect 3096 14909 3124 14910
rect 3096 14883 3097 14909
rect 3097 14883 3123 14909
rect 3123 14883 3124 14909
rect 3096 14882 3124 14883
rect 3148 14909 3176 14910
rect 3148 14883 3149 14909
rect 3149 14883 3175 14909
rect 3175 14883 3176 14909
rect 3148 14882 3176 14883
rect 20888 14909 20916 14910
rect 20888 14883 20889 14909
rect 20889 14883 20915 14909
rect 20915 14883 20916 14909
rect 20888 14882 20916 14883
rect 20940 14909 20968 14910
rect 20940 14883 20941 14909
rect 20941 14883 20967 14909
rect 20967 14883 20968 14909
rect 20940 14882 20968 14883
rect 20992 14909 21020 14910
rect 20992 14883 20993 14909
rect 20993 14883 21019 14909
rect 21019 14883 21020 14909
rect 20992 14882 21020 14883
rect 21044 14909 21072 14910
rect 21044 14883 21045 14909
rect 21045 14883 21071 14909
rect 21071 14883 21072 14909
rect 21044 14882 21072 14883
rect 21096 14909 21124 14910
rect 21096 14883 21097 14909
rect 21097 14883 21123 14909
rect 21123 14883 21124 14909
rect 21096 14882 21124 14883
rect 21148 14909 21176 14910
rect 21148 14883 21149 14909
rect 21149 14883 21175 14909
rect 21175 14883 21176 14909
rect 21148 14882 21176 14883
rect 1028 14517 1056 14518
rect 1028 14491 1029 14517
rect 1029 14491 1055 14517
rect 1055 14491 1056 14517
rect 1028 14490 1056 14491
rect 1080 14517 1108 14518
rect 1080 14491 1081 14517
rect 1081 14491 1107 14517
rect 1107 14491 1108 14517
rect 1080 14490 1108 14491
rect 1132 14517 1160 14518
rect 1132 14491 1133 14517
rect 1133 14491 1159 14517
rect 1159 14491 1160 14517
rect 1132 14490 1160 14491
rect 1184 14517 1212 14518
rect 1184 14491 1185 14517
rect 1185 14491 1211 14517
rect 1211 14491 1212 14517
rect 1184 14490 1212 14491
rect 1236 14517 1264 14518
rect 1236 14491 1237 14517
rect 1237 14491 1263 14517
rect 1263 14491 1264 14517
rect 1236 14490 1264 14491
rect 1288 14517 1316 14518
rect 1288 14491 1289 14517
rect 1289 14491 1315 14517
rect 1315 14491 1316 14517
rect 1288 14490 1316 14491
rect 19028 14517 19056 14518
rect 19028 14491 19029 14517
rect 19029 14491 19055 14517
rect 19055 14491 19056 14517
rect 19028 14490 19056 14491
rect 19080 14517 19108 14518
rect 19080 14491 19081 14517
rect 19081 14491 19107 14517
rect 19107 14491 19108 14517
rect 19080 14490 19108 14491
rect 19132 14517 19160 14518
rect 19132 14491 19133 14517
rect 19133 14491 19159 14517
rect 19159 14491 19160 14517
rect 19132 14490 19160 14491
rect 19184 14517 19212 14518
rect 19184 14491 19185 14517
rect 19185 14491 19211 14517
rect 19211 14491 19212 14517
rect 19184 14490 19212 14491
rect 19236 14517 19264 14518
rect 19236 14491 19237 14517
rect 19237 14491 19263 14517
rect 19263 14491 19264 14517
rect 19236 14490 19264 14491
rect 19288 14517 19316 14518
rect 19288 14491 19289 14517
rect 19289 14491 19315 14517
rect 19315 14491 19316 14517
rect 19288 14490 19316 14491
rect 2888 14125 2916 14126
rect 2888 14099 2889 14125
rect 2889 14099 2915 14125
rect 2915 14099 2916 14125
rect 2888 14098 2916 14099
rect 2940 14125 2968 14126
rect 2940 14099 2941 14125
rect 2941 14099 2967 14125
rect 2967 14099 2968 14125
rect 2940 14098 2968 14099
rect 2992 14125 3020 14126
rect 2992 14099 2993 14125
rect 2993 14099 3019 14125
rect 3019 14099 3020 14125
rect 2992 14098 3020 14099
rect 3044 14125 3072 14126
rect 3044 14099 3045 14125
rect 3045 14099 3071 14125
rect 3071 14099 3072 14125
rect 3044 14098 3072 14099
rect 3096 14125 3124 14126
rect 3096 14099 3097 14125
rect 3097 14099 3123 14125
rect 3123 14099 3124 14125
rect 3096 14098 3124 14099
rect 3148 14125 3176 14126
rect 3148 14099 3149 14125
rect 3149 14099 3175 14125
rect 3175 14099 3176 14125
rect 3148 14098 3176 14099
rect 20888 14125 20916 14126
rect 20888 14099 20889 14125
rect 20889 14099 20915 14125
rect 20915 14099 20916 14125
rect 20888 14098 20916 14099
rect 20940 14125 20968 14126
rect 20940 14099 20941 14125
rect 20941 14099 20967 14125
rect 20967 14099 20968 14125
rect 20940 14098 20968 14099
rect 20992 14125 21020 14126
rect 20992 14099 20993 14125
rect 20993 14099 21019 14125
rect 21019 14099 21020 14125
rect 20992 14098 21020 14099
rect 21044 14125 21072 14126
rect 21044 14099 21045 14125
rect 21045 14099 21071 14125
rect 21071 14099 21072 14125
rect 21044 14098 21072 14099
rect 21096 14125 21124 14126
rect 21096 14099 21097 14125
rect 21097 14099 21123 14125
rect 21123 14099 21124 14125
rect 21096 14098 21124 14099
rect 21148 14125 21176 14126
rect 21148 14099 21149 14125
rect 21149 14099 21175 14125
rect 21175 14099 21176 14125
rect 21148 14098 21176 14099
rect 1028 13733 1056 13734
rect 1028 13707 1029 13733
rect 1029 13707 1055 13733
rect 1055 13707 1056 13733
rect 1028 13706 1056 13707
rect 1080 13733 1108 13734
rect 1080 13707 1081 13733
rect 1081 13707 1107 13733
rect 1107 13707 1108 13733
rect 1080 13706 1108 13707
rect 1132 13733 1160 13734
rect 1132 13707 1133 13733
rect 1133 13707 1159 13733
rect 1159 13707 1160 13733
rect 1132 13706 1160 13707
rect 1184 13733 1212 13734
rect 1184 13707 1185 13733
rect 1185 13707 1211 13733
rect 1211 13707 1212 13733
rect 1184 13706 1212 13707
rect 1236 13733 1264 13734
rect 1236 13707 1237 13733
rect 1237 13707 1263 13733
rect 1263 13707 1264 13733
rect 1236 13706 1264 13707
rect 1288 13733 1316 13734
rect 1288 13707 1289 13733
rect 1289 13707 1315 13733
rect 1315 13707 1316 13733
rect 1288 13706 1316 13707
rect 19028 13733 19056 13734
rect 19028 13707 19029 13733
rect 19029 13707 19055 13733
rect 19055 13707 19056 13733
rect 19028 13706 19056 13707
rect 19080 13733 19108 13734
rect 19080 13707 19081 13733
rect 19081 13707 19107 13733
rect 19107 13707 19108 13733
rect 19080 13706 19108 13707
rect 19132 13733 19160 13734
rect 19132 13707 19133 13733
rect 19133 13707 19159 13733
rect 19159 13707 19160 13733
rect 19132 13706 19160 13707
rect 19184 13733 19212 13734
rect 19184 13707 19185 13733
rect 19185 13707 19211 13733
rect 19211 13707 19212 13733
rect 19184 13706 19212 13707
rect 19236 13733 19264 13734
rect 19236 13707 19237 13733
rect 19237 13707 19263 13733
rect 19263 13707 19264 13733
rect 19236 13706 19264 13707
rect 19288 13733 19316 13734
rect 19288 13707 19289 13733
rect 19289 13707 19315 13733
rect 19315 13707 19316 13733
rect 19288 13706 19316 13707
rect 2888 13341 2916 13342
rect 2888 13315 2889 13341
rect 2889 13315 2915 13341
rect 2915 13315 2916 13341
rect 2888 13314 2916 13315
rect 2940 13341 2968 13342
rect 2940 13315 2941 13341
rect 2941 13315 2967 13341
rect 2967 13315 2968 13341
rect 2940 13314 2968 13315
rect 2992 13341 3020 13342
rect 2992 13315 2993 13341
rect 2993 13315 3019 13341
rect 3019 13315 3020 13341
rect 2992 13314 3020 13315
rect 3044 13341 3072 13342
rect 3044 13315 3045 13341
rect 3045 13315 3071 13341
rect 3071 13315 3072 13341
rect 3044 13314 3072 13315
rect 3096 13341 3124 13342
rect 3096 13315 3097 13341
rect 3097 13315 3123 13341
rect 3123 13315 3124 13341
rect 3096 13314 3124 13315
rect 3148 13341 3176 13342
rect 3148 13315 3149 13341
rect 3149 13315 3175 13341
rect 3175 13315 3176 13341
rect 3148 13314 3176 13315
rect 20888 13341 20916 13342
rect 20888 13315 20889 13341
rect 20889 13315 20915 13341
rect 20915 13315 20916 13341
rect 20888 13314 20916 13315
rect 20940 13341 20968 13342
rect 20940 13315 20941 13341
rect 20941 13315 20967 13341
rect 20967 13315 20968 13341
rect 20940 13314 20968 13315
rect 20992 13341 21020 13342
rect 20992 13315 20993 13341
rect 20993 13315 21019 13341
rect 21019 13315 21020 13341
rect 20992 13314 21020 13315
rect 21044 13341 21072 13342
rect 21044 13315 21045 13341
rect 21045 13315 21071 13341
rect 21071 13315 21072 13341
rect 21044 13314 21072 13315
rect 21096 13341 21124 13342
rect 21096 13315 21097 13341
rect 21097 13315 21123 13341
rect 21123 13315 21124 13341
rect 21096 13314 21124 13315
rect 21148 13341 21176 13342
rect 21148 13315 21149 13341
rect 21149 13315 21175 13341
rect 21175 13315 21176 13341
rect 21148 13314 21176 13315
rect 1028 12949 1056 12950
rect 1028 12923 1029 12949
rect 1029 12923 1055 12949
rect 1055 12923 1056 12949
rect 1028 12922 1056 12923
rect 1080 12949 1108 12950
rect 1080 12923 1081 12949
rect 1081 12923 1107 12949
rect 1107 12923 1108 12949
rect 1080 12922 1108 12923
rect 1132 12949 1160 12950
rect 1132 12923 1133 12949
rect 1133 12923 1159 12949
rect 1159 12923 1160 12949
rect 1132 12922 1160 12923
rect 1184 12949 1212 12950
rect 1184 12923 1185 12949
rect 1185 12923 1211 12949
rect 1211 12923 1212 12949
rect 1184 12922 1212 12923
rect 1236 12949 1264 12950
rect 1236 12923 1237 12949
rect 1237 12923 1263 12949
rect 1263 12923 1264 12949
rect 1236 12922 1264 12923
rect 1288 12949 1316 12950
rect 1288 12923 1289 12949
rect 1289 12923 1315 12949
rect 1315 12923 1316 12949
rect 1288 12922 1316 12923
rect 19028 12949 19056 12950
rect 19028 12923 19029 12949
rect 19029 12923 19055 12949
rect 19055 12923 19056 12949
rect 19028 12922 19056 12923
rect 19080 12949 19108 12950
rect 19080 12923 19081 12949
rect 19081 12923 19107 12949
rect 19107 12923 19108 12949
rect 19080 12922 19108 12923
rect 19132 12949 19160 12950
rect 19132 12923 19133 12949
rect 19133 12923 19159 12949
rect 19159 12923 19160 12949
rect 19132 12922 19160 12923
rect 19184 12949 19212 12950
rect 19184 12923 19185 12949
rect 19185 12923 19211 12949
rect 19211 12923 19212 12949
rect 19184 12922 19212 12923
rect 19236 12949 19264 12950
rect 19236 12923 19237 12949
rect 19237 12923 19263 12949
rect 19263 12923 19264 12949
rect 19236 12922 19264 12923
rect 19288 12949 19316 12950
rect 19288 12923 19289 12949
rect 19289 12923 19315 12949
rect 19315 12923 19316 12949
rect 19288 12922 19316 12923
rect 910 12502 938 12530
rect 2888 12557 2916 12558
rect 2888 12531 2889 12557
rect 2889 12531 2915 12557
rect 2915 12531 2916 12557
rect 2888 12530 2916 12531
rect 2940 12557 2968 12558
rect 2940 12531 2941 12557
rect 2941 12531 2967 12557
rect 2967 12531 2968 12557
rect 2940 12530 2968 12531
rect 2992 12557 3020 12558
rect 2992 12531 2993 12557
rect 2993 12531 3019 12557
rect 3019 12531 3020 12557
rect 2992 12530 3020 12531
rect 3044 12557 3072 12558
rect 3044 12531 3045 12557
rect 3045 12531 3071 12557
rect 3071 12531 3072 12557
rect 3044 12530 3072 12531
rect 3096 12557 3124 12558
rect 3096 12531 3097 12557
rect 3097 12531 3123 12557
rect 3123 12531 3124 12557
rect 3096 12530 3124 12531
rect 3148 12557 3176 12558
rect 3148 12531 3149 12557
rect 3149 12531 3175 12557
rect 3175 12531 3176 12557
rect 3148 12530 3176 12531
rect 20888 12557 20916 12558
rect 20888 12531 20889 12557
rect 20889 12531 20915 12557
rect 20915 12531 20916 12557
rect 20888 12530 20916 12531
rect 20940 12557 20968 12558
rect 20940 12531 20941 12557
rect 20941 12531 20967 12557
rect 20967 12531 20968 12557
rect 20940 12530 20968 12531
rect 20992 12557 21020 12558
rect 20992 12531 20993 12557
rect 20993 12531 21019 12557
rect 21019 12531 21020 12557
rect 20992 12530 21020 12531
rect 21044 12557 21072 12558
rect 21044 12531 21045 12557
rect 21045 12531 21071 12557
rect 21071 12531 21072 12557
rect 21044 12530 21072 12531
rect 21096 12557 21124 12558
rect 21096 12531 21097 12557
rect 21097 12531 21123 12557
rect 21123 12531 21124 12557
rect 21096 12530 21124 12531
rect 21148 12557 21176 12558
rect 21148 12531 21149 12557
rect 21149 12531 21175 12557
rect 21175 12531 21176 12557
rect 21148 12530 21176 12531
rect 22246 12446 22274 12474
rect 1028 12165 1056 12166
rect 1028 12139 1029 12165
rect 1029 12139 1055 12165
rect 1055 12139 1056 12165
rect 1028 12138 1056 12139
rect 1080 12165 1108 12166
rect 1080 12139 1081 12165
rect 1081 12139 1107 12165
rect 1107 12139 1108 12165
rect 1080 12138 1108 12139
rect 1132 12165 1160 12166
rect 1132 12139 1133 12165
rect 1133 12139 1159 12165
rect 1159 12139 1160 12165
rect 1132 12138 1160 12139
rect 1184 12165 1212 12166
rect 1184 12139 1185 12165
rect 1185 12139 1211 12165
rect 1211 12139 1212 12165
rect 1184 12138 1212 12139
rect 1236 12165 1264 12166
rect 1236 12139 1237 12165
rect 1237 12139 1263 12165
rect 1263 12139 1264 12165
rect 1236 12138 1264 12139
rect 1288 12165 1316 12166
rect 1288 12139 1289 12165
rect 1289 12139 1315 12165
rect 1315 12139 1316 12165
rect 1288 12138 1316 12139
rect 19028 12165 19056 12166
rect 19028 12139 19029 12165
rect 19029 12139 19055 12165
rect 19055 12139 19056 12165
rect 19028 12138 19056 12139
rect 19080 12165 19108 12166
rect 19080 12139 19081 12165
rect 19081 12139 19107 12165
rect 19107 12139 19108 12165
rect 19080 12138 19108 12139
rect 19132 12165 19160 12166
rect 19132 12139 19133 12165
rect 19133 12139 19159 12165
rect 19159 12139 19160 12165
rect 19132 12138 19160 12139
rect 19184 12165 19212 12166
rect 19184 12139 19185 12165
rect 19185 12139 19211 12165
rect 19211 12139 19212 12165
rect 19184 12138 19212 12139
rect 19236 12165 19264 12166
rect 19236 12139 19237 12165
rect 19237 12139 19263 12165
rect 19263 12139 19264 12165
rect 19236 12138 19264 12139
rect 19288 12165 19316 12166
rect 19288 12139 19289 12165
rect 19289 12139 19315 12165
rect 19315 12139 19316 12165
rect 19288 12138 19316 12139
rect 2888 11773 2916 11774
rect 2888 11747 2889 11773
rect 2889 11747 2915 11773
rect 2915 11747 2916 11773
rect 2888 11746 2916 11747
rect 2940 11773 2968 11774
rect 2940 11747 2941 11773
rect 2941 11747 2967 11773
rect 2967 11747 2968 11773
rect 2940 11746 2968 11747
rect 2992 11773 3020 11774
rect 2992 11747 2993 11773
rect 2993 11747 3019 11773
rect 3019 11747 3020 11773
rect 2992 11746 3020 11747
rect 3044 11773 3072 11774
rect 3044 11747 3045 11773
rect 3045 11747 3071 11773
rect 3071 11747 3072 11773
rect 3044 11746 3072 11747
rect 3096 11773 3124 11774
rect 3096 11747 3097 11773
rect 3097 11747 3123 11773
rect 3123 11747 3124 11773
rect 3096 11746 3124 11747
rect 3148 11773 3176 11774
rect 3148 11747 3149 11773
rect 3149 11747 3175 11773
rect 3175 11747 3176 11773
rect 3148 11746 3176 11747
rect 20888 11773 20916 11774
rect 20888 11747 20889 11773
rect 20889 11747 20915 11773
rect 20915 11747 20916 11773
rect 20888 11746 20916 11747
rect 20940 11773 20968 11774
rect 20940 11747 20941 11773
rect 20941 11747 20967 11773
rect 20967 11747 20968 11773
rect 20940 11746 20968 11747
rect 20992 11773 21020 11774
rect 20992 11747 20993 11773
rect 20993 11747 21019 11773
rect 21019 11747 21020 11773
rect 20992 11746 21020 11747
rect 21044 11773 21072 11774
rect 21044 11747 21045 11773
rect 21045 11747 21071 11773
rect 21071 11747 21072 11773
rect 21044 11746 21072 11747
rect 21096 11773 21124 11774
rect 21096 11747 21097 11773
rect 21097 11747 21123 11773
rect 21123 11747 21124 11773
rect 21096 11746 21124 11747
rect 21148 11773 21176 11774
rect 21148 11747 21149 11773
rect 21149 11747 21175 11773
rect 21175 11747 21176 11773
rect 21148 11746 21176 11747
rect 1028 11381 1056 11382
rect 1028 11355 1029 11381
rect 1029 11355 1055 11381
rect 1055 11355 1056 11381
rect 1028 11354 1056 11355
rect 1080 11381 1108 11382
rect 1080 11355 1081 11381
rect 1081 11355 1107 11381
rect 1107 11355 1108 11381
rect 1080 11354 1108 11355
rect 1132 11381 1160 11382
rect 1132 11355 1133 11381
rect 1133 11355 1159 11381
rect 1159 11355 1160 11381
rect 1132 11354 1160 11355
rect 1184 11381 1212 11382
rect 1184 11355 1185 11381
rect 1185 11355 1211 11381
rect 1211 11355 1212 11381
rect 1184 11354 1212 11355
rect 1236 11381 1264 11382
rect 1236 11355 1237 11381
rect 1237 11355 1263 11381
rect 1263 11355 1264 11381
rect 1236 11354 1264 11355
rect 1288 11381 1316 11382
rect 1288 11355 1289 11381
rect 1289 11355 1315 11381
rect 1315 11355 1316 11381
rect 1288 11354 1316 11355
rect 19028 11381 19056 11382
rect 19028 11355 19029 11381
rect 19029 11355 19055 11381
rect 19055 11355 19056 11381
rect 19028 11354 19056 11355
rect 19080 11381 19108 11382
rect 19080 11355 19081 11381
rect 19081 11355 19107 11381
rect 19107 11355 19108 11381
rect 19080 11354 19108 11355
rect 19132 11381 19160 11382
rect 19132 11355 19133 11381
rect 19133 11355 19159 11381
rect 19159 11355 19160 11381
rect 19132 11354 19160 11355
rect 19184 11381 19212 11382
rect 19184 11355 19185 11381
rect 19185 11355 19211 11381
rect 19211 11355 19212 11381
rect 19184 11354 19212 11355
rect 19236 11381 19264 11382
rect 19236 11355 19237 11381
rect 19237 11355 19263 11381
rect 19263 11355 19264 11381
rect 19236 11354 19264 11355
rect 19288 11381 19316 11382
rect 19288 11355 19289 11381
rect 19289 11355 19315 11381
rect 19315 11355 19316 11381
rect 19288 11354 19316 11355
rect 2888 10989 2916 10990
rect 2888 10963 2889 10989
rect 2889 10963 2915 10989
rect 2915 10963 2916 10989
rect 2888 10962 2916 10963
rect 2940 10989 2968 10990
rect 2940 10963 2941 10989
rect 2941 10963 2967 10989
rect 2967 10963 2968 10989
rect 2940 10962 2968 10963
rect 2992 10989 3020 10990
rect 2992 10963 2993 10989
rect 2993 10963 3019 10989
rect 3019 10963 3020 10989
rect 2992 10962 3020 10963
rect 3044 10989 3072 10990
rect 3044 10963 3045 10989
rect 3045 10963 3071 10989
rect 3071 10963 3072 10989
rect 3044 10962 3072 10963
rect 3096 10989 3124 10990
rect 3096 10963 3097 10989
rect 3097 10963 3123 10989
rect 3123 10963 3124 10989
rect 3096 10962 3124 10963
rect 3148 10989 3176 10990
rect 3148 10963 3149 10989
rect 3149 10963 3175 10989
rect 3175 10963 3176 10989
rect 3148 10962 3176 10963
rect 20888 10989 20916 10990
rect 20888 10963 20889 10989
rect 20889 10963 20915 10989
rect 20915 10963 20916 10989
rect 20888 10962 20916 10963
rect 20940 10989 20968 10990
rect 20940 10963 20941 10989
rect 20941 10963 20967 10989
rect 20967 10963 20968 10989
rect 20940 10962 20968 10963
rect 20992 10989 21020 10990
rect 20992 10963 20993 10989
rect 20993 10963 21019 10989
rect 21019 10963 21020 10989
rect 20992 10962 21020 10963
rect 21044 10989 21072 10990
rect 21044 10963 21045 10989
rect 21045 10963 21071 10989
rect 21071 10963 21072 10989
rect 21044 10962 21072 10963
rect 21096 10989 21124 10990
rect 21096 10963 21097 10989
rect 21097 10963 21123 10989
rect 21123 10963 21124 10989
rect 21096 10962 21124 10963
rect 21148 10989 21176 10990
rect 21148 10963 21149 10989
rect 21149 10963 21175 10989
rect 21175 10963 21176 10989
rect 21148 10962 21176 10963
rect 1028 10597 1056 10598
rect 1028 10571 1029 10597
rect 1029 10571 1055 10597
rect 1055 10571 1056 10597
rect 1028 10570 1056 10571
rect 1080 10597 1108 10598
rect 1080 10571 1081 10597
rect 1081 10571 1107 10597
rect 1107 10571 1108 10597
rect 1080 10570 1108 10571
rect 1132 10597 1160 10598
rect 1132 10571 1133 10597
rect 1133 10571 1159 10597
rect 1159 10571 1160 10597
rect 1132 10570 1160 10571
rect 1184 10597 1212 10598
rect 1184 10571 1185 10597
rect 1185 10571 1211 10597
rect 1211 10571 1212 10597
rect 1184 10570 1212 10571
rect 1236 10597 1264 10598
rect 1236 10571 1237 10597
rect 1237 10571 1263 10597
rect 1263 10571 1264 10597
rect 1236 10570 1264 10571
rect 1288 10597 1316 10598
rect 1288 10571 1289 10597
rect 1289 10571 1315 10597
rect 1315 10571 1316 10597
rect 1288 10570 1316 10571
rect 19028 10597 19056 10598
rect 19028 10571 19029 10597
rect 19029 10571 19055 10597
rect 19055 10571 19056 10597
rect 19028 10570 19056 10571
rect 19080 10597 19108 10598
rect 19080 10571 19081 10597
rect 19081 10571 19107 10597
rect 19107 10571 19108 10597
rect 19080 10570 19108 10571
rect 19132 10597 19160 10598
rect 19132 10571 19133 10597
rect 19133 10571 19159 10597
rect 19159 10571 19160 10597
rect 19132 10570 19160 10571
rect 19184 10597 19212 10598
rect 19184 10571 19185 10597
rect 19185 10571 19211 10597
rect 19211 10571 19212 10597
rect 19184 10570 19212 10571
rect 19236 10597 19264 10598
rect 19236 10571 19237 10597
rect 19237 10571 19263 10597
rect 19263 10571 19264 10597
rect 19236 10570 19264 10571
rect 19288 10597 19316 10598
rect 19288 10571 19289 10597
rect 19289 10571 19315 10597
rect 19315 10571 19316 10597
rect 19288 10570 19316 10571
rect 2888 10205 2916 10206
rect 2888 10179 2889 10205
rect 2889 10179 2915 10205
rect 2915 10179 2916 10205
rect 2888 10178 2916 10179
rect 2940 10205 2968 10206
rect 2940 10179 2941 10205
rect 2941 10179 2967 10205
rect 2967 10179 2968 10205
rect 2940 10178 2968 10179
rect 2992 10205 3020 10206
rect 2992 10179 2993 10205
rect 2993 10179 3019 10205
rect 3019 10179 3020 10205
rect 2992 10178 3020 10179
rect 3044 10205 3072 10206
rect 3044 10179 3045 10205
rect 3045 10179 3071 10205
rect 3071 10179 3072 10205
rect 3044 10178 3072 10179
rect 3096 10205 3124 10206
rect 3096 10179 3097 10205
rect 3097 10179 3123 10205
rect 3123 10179 3124 10205
rect 3096 10178 3124 10179
rect 3148 10205 3176 10206
rect 3148 10179 3149 10205
rect 3149 10179 3175 10205
rect 3175 10179 3176 10205
rect 3148 10178 3176 10179
rect 20888 10205 20916 10206
rect 20888 10179 20889 10205
rect 20889 10179 20915 10205
rect 20915 10179 20916 10205
rect 20888 10178 20916 10179
rect 20940 10205 20968 10206
rect 20940 10179 20941 10205
rect 20941 10179 20967 10205
rect 20967 10179 20968 10205
rect 20940 10178 20968 10179
rect 20992 10205 21020 10206
rect 20992 10179 20993 10205
rect 20993 10179 21019 10205
rect 21019 10179 21020 10205
rect 20992 10178 21020 10179
rect 21044 10205 21072 10206
rect 21044 10179 21045 10205
rect 21045 10179 21071 10205
rect 21071 10179 21072 10205
rect 21044 10178 21072 10179
rect 21096 10205 21124 10206
rect 21096 10179 21097 10205
rect 21097 10179 21123 10205
rect 21123 10179 21124 10205
rect 21096 10178 21124 10179
rect 21148 10205 21176 10206
rect 21148 10179 21149 10205
rect 21149 10179 21175 10205
rect 21175 10179 21176 10205
rect 21148 10178 21176 10179
rect 1028 9813 1056 9814
rect 1028 9787 1029 9813
rect 1029 9787 1055 9813
rect 1055 9787 1056 9813
rect 1028 9786 1056 9787
rect 1080 9813 1108 9814
rect 1080 9787 1081 9813
rect 1081 9787 1107 9813
rect 1107 9787 1108 9813
rect 1080 9786 1108 9787
rect 1132 9813 1160 9814
rect 1132 9787 1133 9813
rect 1133 9787 1159 9813
rect 1159 9787 1160 9813
rect 1132 9786 1160 9787
rect 1184 9813 1212 9814
rect 1184 9787 1185 9813
rect 1185 9787 1211 9813
rect 1211 9787 1212 9813
rect 1184 9786 1212 9787
rect 1236 9813 1264 9814
rect 1236 9787 1237 9813
rect 1237 9787 1263 9813
rect 1263 9787 1264 9813
rect 1236 9786 1264 9787
rect 1288 9813 1316 9814
rect 1288 9787 1289 9813
rect 1289 9787 1315 9813
rect 1315 9787 1316 9813
rect 1288 9786 1316 9787
rect 19028 9813 19056 9814
rect 19028 9787 19029 9813
rect 19029 9787 19055 9813
rect 19055 9787 19056 9813
rect 19028 9786 19056 9787
rect 19080 9813 19108 9814
rect 19080 9787 19081 9813
rect 19081 9787 19107 9813
rect 19107 9787 19108 9813
rect 19080 9786 19108 9787
rect 19132 9813 19160 9814
rect 19132 9787 19133 9813
rect 19133 9787 19159 9813
rect 19159 9787 19160 9813
rect 19132 9786 19160 9787
rect 19184 9813 19212 9814
rect 19184 9787 19185 9813
rect 19185 9787 19211 9813
rect 19211 9787 19212 9813
rect 19184 9786 19212 9787
rect 19236 9813 19264 9814
rect 19236 9787 19237 9813
rect 19237 9787 19263 9813
rect 19263 9787 19264 9813
rect 19236 9786 19264 9787
rect 19288 9813 19316 9814
rect 19288 9787 19289 9813
rect 19289 9787 19315 9813
rect 19315 9787 19316 9813
rect 19288 9786 19316 9787
rect 2888 9421 2916 9422
rect 2888 9395 2889 9421
rect 2889 9395 2915 9421
rect 2915 9395 2916 9421
rect 2888 9394 2916 9395
rect 2940 9421 2968 9422
rect 2940 9395 2941 9421
rect 2941 9395 2967 9421
rect 2967 9395 2968 9421
rect 2940 9394 2968 9395
rect 2992 9421 3020 9422
rect 2992 9395 2993 9421
rect 2993 9395 3019 9421
rect 3019 9395 3020 9421
rect 2992 9394 3020 9395
rect 3044 9421 3072 9422
rect 3044 9395 3045 9421
rect 3045 9395 3071 9421
rect 3071 9395 3072 9421
rect 3044 9394 3072 9395
rect 3096 9421 3124 9422
rect 3096 9395 3097 9421
rect 3097 9395 3123 9421
rect 3123 9395 3124 9421
rect 3096 9394 3124 9395
rect 3148 9421 3176 9422
rect 3148 9395 3149 9421
rect 3149 9395 3175 9421
rect 3175 9395 3176 9421
rect 3148 9394 3176 9395
rect 20888 9421 20916 9422
rect 20888 9395 20889 9421
rect 20889 9395 20915 9421
rect 20915 9395 20916 9421
rect 20888 9394 20916 9395
rect 20940 9421 20968 9422
rect 20940 9395 20941 9421
rect 20941 9395 20967 9421
rect 20967 9395 20968 9421
rect 20940 9394 20968 9395
rect 20992 9421 21020 9422
rect 20992 9395 20993 9421
rect 20993 9395 21019 9421
rect 21019 9395 21020 9421
rect 20992 9394 21020 9395
rect 21044 9421 21072 9422
rect 21044 9395 21045 9421
rect 21045 9395 21071 9421
rect 21071 9395 21072 9421
rect 21044 9394 21072 9395
rect 21096 9421 21124 9422
rect 21096 9395 21097 9421
rect 21097 9395 21123 9421
rect 21123 9395 21124 9421
rect 21096 9394 21124 9395
rect 21148 9421 21176 9422
rect 21148 9395 21149 9421
rect 21149 9395 21175 9421
rect 21175 9395 21176 9421
rect 21148 9394 21176 9395
rect 1028 9029 1056 9030
rect 1028 9003 1029 9029
rect 1029 9003 1055 9029
rect 1055 9003 1056 9029
rect 1028 9002 1056 9003
rect 1080 9029 1108 9030
rect 1080 9003 1081 9029
rect 1081 9003 1107 9029
rect 1107 9003 1108 9029
rect 1080 9002 1108 9003
rect 1132 9029 1160 9030
rect 1132 9003 1133 9029
rect 1133 9003 1159 9029
rect 1159 9003 1160 9029
rect 1132 9002 1160 9003
rect 1184 9029 1212 9030
rect 1184 9003 1185 9029
rect 1185 9003 1211 9029
rect 1211 9003 1212 9029
rect 1184 9002 1212 9003
rect 1236 9029 1264 9030
rect 1236 9003 1237 9029
rect 1237 9003 1263 9029
rect 1263 9003 1264 9029
rect 1236 9002 1264 9003
rect 1288 9029 1316 9030
rect 1288 9003 1289 9029
rect 1289 9003 1315 9029
rect 1315 9003 1316 9029
rect 1288 9002 1316 9003
rect 19028 9029 19056 9030
rect 19028 9003 19029 9029
rect 19029 9003 19055 9029
rect 19055 9003 19056 9029
rect 19028 9002 19056 9003
rect 19080 9029 19108 9030
rect 19080 9003 19081 9029
rect 19081 9003 19107 9029
rect 19107 9003 19108 9029
rect 19080 9002 19108 9003
rect 19132 9029 19160 9030
rect 19132 9003 19133 9029
rect 19133 9003 19159 9029
rect 19159 9003 19160 9029
rect 19132 9002 19160 9003
rect 19184 9029 19212 9030
rect 19184 9003 19185 9029
rect 19185 9003 19211 9029
rect 19211 9003 19212 9029
rect 19184 9002 19212 9003
rect 19236 9029 19264 9030
rect 19236 9003 19237 9029
rect 19237 9003 19263 9029
rect 19263 9003 19264 9029
rect 19236 9002 19264 9003
rect 19288 9029 19316 9030
rect 19288 9003 19289 9029
rect 19289 9003 19315 9029
rect 19315 9003 19316 9029
rect 19288 9002 19316 9003
rect 2888 8637 2916 8638
rect 2888 8611 2889 8637
rect 2889 8611 2915 8637
rect 2915 8611 2916 8637
rect 2888 8610 2916 8611
rect 2940 8637 2968 8638
rect 2940 8611 2941 8637
rect 2941 8611 2967 8637
rect 2967 8611 2968 8637
rect 2940 8610 2968 8611
rect 2992 8637 3020 8638
rect 2992 8611 2993 8637
rect 2993 8611 3019 8637
rect 3019 8611 3020 8637
rect 2992 8610 3020 8611
rect 3044 8637 3072 8638
rect 3044 8611 3045 8637
rect 3045 8611 3071 8637
rect 3071 8611 3072 8637
rect 3044 8610 3072 8611
rect 3096 8637 3124 8638
rect 3096 8611 3097 8637
rect 3097 8611 3123 8637
rect 3123 8611 3124 8637
rect 3096 8610 3124 8611
rect 3148 8637 3176 8638
rect 3148 8611 3149 8637
rect 3149 8611 3175 8637
rect 3175 8611 3176 8637
rect 3148 8610 3176 8611
rect 20888 8637 20916 8638
rect 20888 8611 20889 8637
rect 20889 8611 20915 8637
rect 20915 8611 20916 8637
rect 20888 8610 20916 8611
rect 20940 8637 20968 8638
rect 20940 8611 20941 8637
rect 20941 8611 20967 8637
rect 20967 8611 20968 8637
rect 20940 8610 20968 8611
rect 20992 8637 21020 8638
rect 20992 8611 20993 8637
rect 20993 8611 21019 8637
rect 21019 8611 21020 8637
rect 20992 8610 21020 8611
rect 21044 8637 21072 8638
rect 21044 8611 21045 8637
rect 21045 8611 21071 8637
rect 21071 8611 21072 8637
rect 21044 8610 21072 8611
rect 21096 8637 21124 8638
rect 21096 8611 21097 8637
rect 21097 8611 21123 8637
rect 21123 8611 21124 8637
rect 21096 8610 21124 8611
rect 21148 8637 21176 8638
rect 21148 8611 21149 8637
rect 21149 8611 21175 8637
rect 21175 8611 21176 8637
rect 21148 8610 21176 8611
rect 1028 8245 1056 8246
rect 1028 8219 1029 8245
rect 1029 8219 1055 8245
rect 1055 8219 1056 8245
rect 1028 8218 1056 8219
rect 1080 8245 1108 8246
rect 1080 8219 1081 8245
rect 1081 8219 1107 8245
rect 1107 8219 1108 8245
rect 1080 8218 1108 8219
rect 1132 8245 1160 8246
rect 1132 8219 1133 8245
rect 1133 8219 1159 8245
rect 1159 8219 1160 8245
rect 1132 8218 1160 8219
rect 1184 8245 1212 8246
rect 1184 8219 1185 8245
rect 1185 8219 1211 8245
rect 1211 8219 1212 8245
rect 1184 8218 1212 8219
rect 1236 8245 1264 8246
rect 1236 8219 1237 8245
rect 1237 8219 1263 8245
rect 1263 8219 1264 8245
rect 1236 8218 1264 8219
rect 1288 8245 1316 8246
rect 1288 8219 1289 8245
rect 1289 8219 1315 8245
rect 1315 8219 1316 8245
rect 1288 8218 1316 8219
rect 19028 8245 19056 8246
rect 19028 8219 19029 8245
rect 19029 8219 19055 8245
rect 19055 8219 19056 8245
rect 19028 8218 19056 8219
rect 19080 8245 19108 8246
rect 19080 8219 19081 8245
rect 19081 8219 19107 8245
rect 19107 8219 19108 8245
rect 19080 8218 19108 8219
rect 19132 8245 19160 8246
rect 19132 8219 19133 8245
rect 19133 8219 19159 8245
rect 19159 8219 19160 8245
rect 19132 8218 19160 8219
rect 19184 8245 19212 8246
rect 19184 8219 19185 8245
rect 19185 8219 19211 8245
rect 19211 8219 19212 8245
rect 19184 8218 19212 8219
rect 19236 8245 19264 8246
rect 19236 8219 19237 8245
rect 19237 8219 19263 8245
rect 19263 8219 19264 8245
rect 19236 8218 19264 8219
rect 19288 8245 19316 8246
rect 19288 8219 19289 8245
rect 19289 8219 19315 8245
rect 19315 8219 19316 8245
rect 19288 8218 19316 8219
rect 2888 7853 2916 7854
rect 2888 7827 2889 7853
rect 2889 7827 2915 7853
rect 2915 7827 2916 7853
rect 2888 7826 2916 7827
rect 2940 7853 2968 7854
rect 2940 7827 2941 7853
rect 2941 7827 2967 7853
rect 2967 7827 2968 7853
rect 2940 7826 2968 7827
rect 2992 7853 3020 7854
rect 2992 7827 2993 7853
rect 2993 7827 3019 7853
rect 3019 7827 3020 7853
rect 2992 7826 3020 7827
rect 3044 7853 3072 7854
rect 3044 7827 3045 7853
rect 3045 7827 3071 7853
rect 3071 7827 3072 7853
rect 3044 7826 3072 7827
rect 3096 7853 3124 7854
rect 3096 7827 3097 7853
rect 3097 7827 3123 7853
rect 3123 7827 3124 7853
rect 3096 7826 3124 7827
rect 3148 7853 3176 7854
rect 3148 7827 3149 7853
rect 3149 7827 3175 7853
rect 3175 7827 3176 7853
rect 3148 7826 3176 7827
rect 20888 7853 20916 7854
rect 20888 7827 20889 7853
rect 20889 7827 20915 7853
rect 20915 7827 20916 7853
rect 20888 7826 20916 7827
rect 20940 7853 20968 7854
rect 20940 7827 20941 7853
rect 20941 7827 20967 7853
rect 20967 7827 20968 7853
rect 20940 7826 20968 7827
rect 20992 7853 21020 7854
rect 20992 7827 20993 7853
rect 20993 7827 21019 7853
rect 21019 7827 21020 7853
rect 20992 7826 21020 7827
rect 21044 7853 21072 7854
rect 21044 7827 21045 7853
rect 21045 7827 21071 7853
rect 21071 7827 21072 7853
rect 21044 7826 21072 7827
rect 21096 7853 21124 7854
rect 21096 7827 21097 7853
rect 21097 7827 21123 7853
rect 21123 7827 21124 7853
rect 21096 7826 21124 7827
rect 21148 7853 21176 7854
rect 21148 7827 21149 7853
rect 21149 7827 21175 7853
rect 21175 7827 21176 7853
rect 21148 7826 21176 7827
rect 1028 7461 1056 7462
rect 1028 7435 1029 7461
rect 1029 7435 1055 7461
rect 1055 7435 1056 7461
rect 1028 7434 1056 7435
rect 1080 7461 1108 7462
rect 1080 7435 1081 7461
rect 1081 7435 1107 7461
rect 1107 7435 1108 7461
rect 1080 7434 1108 7435
rect 1132 7461 1160 7462
rect 1132 7435 1133 7461
rect 1133 7435 1159 7461
rect 1159 7435 1160 7461
rect 1132 7434 1160 7435
rect 1184 7461 1212 7462
rect 1184 7435 1185 7461
rect 1185 7435 1211 7461
rect 1211 7435 1212 7461
rect 1184 7434 1212 7435
rect 1236 7461 1264 7462
rect 1236 7435 1237 7461
rect 1237 7435 1263 7461
rect 1263 7435 1264 7461
rect 1236 7434 1264 7435
rect 1288 7461 1316 7462
rect 1288 7435 1289 7461
rect 1289 7435 1315 7461
rect 1315 7435 1316 7461
rect 1288 7434 1316 7435
rect 19028 7461 19056 7462
rect 19028 7435 19029 7461
rect 19029 7435 19055 7461
rect 19055 7435 19056 7461
rect 19028 7434 19056 7435
rect 19080 7461 19108 7462
rect 19080 7435 19081 7461
rect 19081 7435 19107 7461
rect 19107 7435 19108 7461
rect 19080 7434 19108 7435
rect 19132 7461 19160 7462
rect 19132 7435 19133 7461
rect 19133 7435 19159 7461
rect 19159 7435 19160 7461
rect 19132 7434 19160 7435
rect 19184 7461 19212 7462
rect 19184 7435 19185 7461
rect 19185 7435 19211 7461
rect 19211 7435 19212 7461
rect 19184 7434 19212 7435
rect 19236 7461 19264 7462
rect 19236 7435 19237 7461
rect 19237 7435 19263 7461
rect 19263 7435 19264 7461
rect 19236 7434 19264 7435
rect 19288 7461 19316 7462
rect 19288 7435 19289 7461
rect 19289 7435 19315 7461
rect 19315 7435 19316 7461
rect 19288 7434 19316 7435
rect 2888 7069 2916 7070
rect 2888 7043 2889 7069
rect 2889 7043 2915 7069
rect 2915 7043 2916 7069
rect 2888 7042 2916 7043
rect 2940 7069 2968 7070
rect 2940 7043 2941 7069
rect 2941 7043 2967 7069
rect 2967 7043 2968 7069
rect 2940 7042 2968 7043
rect 2992 7069 3020 7070
rect 2992 7043 2993 7069
rect 2993 7043 3019 7069
rect 3019 7043 3020 7069
rect 2992 7042 3020 7043
rect 3044 7069 3072 7070
rect 3044 7043 3045 7069
rect 3045 7043 3071 7069
rect 3071 7043 3072 7069
rect 3044 7042 3072 7043
rect 3096 7069 3124 7070
rect 3096 7043 3097 7069
rect 3097 7043 3123 7069
rect 3123 7043 3124 7069
rect 3096 7042 3124 7043
rect 3148 7069 3176 7070
rect 3148 7043 3149 7069
rect 3149 7043 3175 7069
rect 3175 7043 3176 7069
rect 3148 7042 3176 7043
rect 20888 7069 20916 7070
rect 20888 7043 20889 7069
rect 20889 7043 20915 7069
rect 20915 7043 20916 7069
rect 20888 7042 20916 7043
rect 20940 7069 20968 7070
rect 20940 7043 20941 7069
rect 20941 7043 20967 7069
rect 20967 7043 20968 7069
rect 20940 7042 20968 7043
rect 20992 7069 21020 7070
rect 20992 7043 20993 7069
rect 20993 7043 21019 7069
rect 21019 7043 21020 7069
rect 20992 7042 21020 7043
rect 21044 7069 21072 7070
rect 21044 7043 21045 7069
rect 21045 7043 21071 7069
rect 21071 7043 21072 7069
rect 21044 7042 21072 7043
rect 21096 7069 21124 7070
rect 21096 7043 21097 7069
rect 21097 7043 21123 7069
rect 21123 7043 21124 7069
rect 21096 7042 21124 7043
rect 21148 7069 21176 7070
rect 21148 7043 21149 7069
rect 21149 7043 21175 7069
rect 21175 7043 21176 7069
rect 21148 7042 21176 7043
rect 1028 6677 1056 6678
rect 1028 6651 1029 6677
rect 1029 6651 1055 6677
rect 1055 6651 1056 6677
rect 1028 6650 1056 6651
rect 1080 6677 1108 6678
rect 1080 6651 1081 6677
rect 1081 6651 1107 6677
rect 1107 6651 1108 6677
rect 1080 6650 1108 6651
rect 1132 6677 1160 6678
rect 1132 6651 1133 6677
rect 1133 6651 1159 6677
rect 1159 6651 1160 6677
rect 1132 6650 1160 6651
rect 1184 6677 1212 6678
rect 1184 6651 1185 6677
rect 1185 6651 1211 6677
rect 1211 6651 1212 6677
rect 1184 6650 1212 6651
rect 1236 6677 1264 6678
rect 1236 6651 1237 6677
rect 1237 6651 1263 6677
rect 1263 6651 1264 6677
rect 1236 6650 1264 6651
rect 1288 6677 1316 6678
rect 1288 6651 1289 6677
rect 1289 6651 1315 6677
rect 1315 6651 1316 6677
rect 1288 6650 1316 6651
rect 19028 6677 19056 6678
rect 19028 6651 19029 6677
rect 19029 6651 19055 6677
rect 19055 6651 19056 6677
rect 19028 6650 19056 6651
rect 19080 6677 19108 6678
rect 19080 6651 19081 6677
rect 19081 6651 19107 6677
rect 19107 6651 19108 6677
rect 19080 6650 19108 6651
rect 19132 6677 19160 6678
rect 19132 6651 19133 6677
rect 19133 6651 19159 6677
rect 19159 6651 19160 6677
rect 19132 6650 19160 6651
rect 19184 6677 19212 6678
rect 19184 6651 19185 6677
rect 19185 6651 19211 6677
rect 19211 6651 19212 6677
rect 19184 6650 19212 6651
rect 19236 6677 19264 6678
rect 19236 6651 19237 6677
rect 19237 6651 19263 6677
rect 19263 6651 19264 6677
rect 19236 6650 19264 6651
rect 19288 6677 19316 6678
rect 19288 6651 19289 6677
rect 19289 6651 19315 6677
rect 19315 6651 19316 6677
rect 19288 6650 19316 6651
rect 2888 6285 2916 6286
rect 2888 6259 2889 6285
rect 2889 6259 2915 6285
rect 2915 6259 2916 6285
rect 2888 6258 2916 6259
rect 2940 6285 2968 6286
rect 2940 6259 2941 6285
rect 2941 6259 2967 6285
rect 2967 6259 2968 6285
rect 2940 6258 2968 6259
rect 2992 6285 3020 6286
rect 2992 6259 2993 6285
rect 2993 6259 3019 6285
rect 3019 6259 3020 6285
rect 2992 6258 3020 6259
rect 3044 6285 3072 6286
rect 3044 6259 3045 6285
rect 3045 6259 3071 6285
rect 3071 6259 3072 6285
rect 3044 6258 3072 6259
rect 3096 6285 3124 6286
rect 3096 6259 3097 6285
rect 3097 6259 3123 6285
rect 3123 6259 3124 6285
rect 3096 6258 3124 6259
rect 3148 6285 3176 6286
rect 3148 6259 3149 6285
rect 3149 6259 3175 6285
rect 3175 6259 3176 6285
rect 3148 6258 3176 6259
rect 20888 6285 20916 6286
rect 20888 6259 20889 6285
rect 20889 6259 20915 6285
rect 20915 6259 20916 6285
rect 20888 6258 20916 6259
rect 20940 6285 20968 6286
rect 20940 6259 20941 6285
rect 20941 6259 20967 6285
rect 20967 6259 20968 6285
rect 20940 6258 20968 6259
rect 20992 6285 21020 6286
rect 20992 6259 20993 6285
rect 20993 6259 21019 6285
rect 21019 6259 21020 6285
rect 20992 6258 21020 6259
rect 21044 6285 21072 6286
rect 21044 6259 21045 6285
rect 21045 6259 21071 6285
rect 21071 6259 21072 6285
rect 21044 6258 21072 6259
rect 21096 6285 21124 6286
rect 21096 6259 21097 6285
rect 21097 6259 21123 6285
rect 21123 6259 21124 6285
rect 21096 6258 21124 6259
rect 21148 6285 21176 6286
rect 21148 6259 21149 6285
rect 21149 6259 21175 6285
rect 21175 6259 21176 6285
rect 21148 6258 21176 6259
rect 14294 6062 14322 6090
rect 12894 6006 12922 6034
rect 1028 5893 1056 5894
rect 1028 5867 1029 5893
rect 1029 5867 1055 5893
rect 1055 5867 1056 5893
rect 1028 5866 1056 5867
rect 1080 5893 1108 5894
rect 1080 5867 1081 5893
rect 1081 5867 1107 5893
rect 1107 5867 1108 5893
rect 1080 5866 1108 5867
rect 1132 5893 1160 5894
rect 1132 5867 1133 5893
rect 1133 5867 1159 5893
rect 1159 5867 1160 5893
rect 1132 5866 1160 5867
rect 1184 5893 1212 5894
rect 1184 5867 1185 5893
rect 1185 5867 1211 5893
rect 1211 5867 1212 5893
rect 1184 5866 1212 5867
rect 1236 5893 1264 5894
rect 1236 5867 1237 5893
rect 1237 5867 1263 5893
rect 1263 5867 1264 5893
rect 1236 5866 1264 5867
rect 1288 5893 1316 5894
rect 1288 5867 1289 5893
rect 1289 5867 1315 5893
rect 1315 5867 1316 5893
rect 1288 5866 1316 5867
rect 2888 5501 2916 5502
rect 2888 5475 2889 5501
rect 2889 5475 2915 5501
rect 2915 5475 2916 5501
rect 2888 5474 2916 5475
rect 2940 5501 2968 5502
rect 2940 5475 2941 5501
rect 2941 5475 2967 5501
rect 2967 5475 2968 5501
rect 2940 5474 2968 5475
rect 2992 5501 3020 5502
rect 2992 5475 2993 5501
rect 2993 5475 3019 5501
rect 3019 5475 3020 5501
rect 2992 5474 3020 5475
rect 3044 5501 3072 5502
rect 3044 5475 3045 5501
rect 3045 5475 3071 5501
rect 3071 5475 3072 5501
rect 3044 5474 3072 5475
rect 3096 5501 3124 5502
rect 3096 5475 3097 5501
rect 3097 5475 3123 5501
rect 3123 5475 3124 5501
rect 3096 5474 3124 5475
rect 3148 5501 3176 5502
rect 3148 5475 3149 5501
rect 3149 5475 3175 5501
rect 3175 5475 3176 5501
rect 3148 5474 3176 5475
rect 12502 5558 12530 5586
rect 13510 6033 13538 6034
rect 13510 6007 13511 6033
rect 13511 6007 13537 6033
rect 13537 6007 13538 6033
rect 13510 6006 13538 6007
rect 13230 5585 13258 5586
rect 13230 5559 13231 5585
rect 13231 5559 13257 5585
rect 13257 5559 13258 5585
rect 13230 5558 13258 5559
rect 6286 5222 6314 5250
rect 1028 5109 1056 5110
rect 1028 5083 1029 5109
rect 1029 5083 1055 5109
rect 1055 5083 1056 5109
rect 1028 5082 1056 5083
rect 1080 5109 1108 5110
rect 1080 5083 1081 5109
rect 1081 5083 1107 5109
rect 1107 5083 1108 5109
rect 1080 5082 1108 5083
rect 1132 5109 1160 5110
rect 1132 5083 1133 5109
rect 1133 5083 1159 5109
rect 1159 5083 1160 5109
rect 1132 5082 1160 5083
rect 1184 5109 1212 5110
rect 1184 5083 1185 5109
rect 1185 5083 1211 5109
rect 1211 5083 1212 5109
rect 1184 5082 1212 5083
rect 1236 5109 1264 5110
rect 1236 5083 1237 5109
rect 1237 5083 1263 5109
rect 1263 5083 1264 5109
rect 1236 5082 1264 5083
rect 1288 5109 1316 5110
rect 1288 5083 1289 5109
rect 1289 5083 1315 5109
rect 1315 5083 1316 5109
rect 1288 5082 1316 5083
rect 2888 4717 2916 4718
rect 2888 4691 2889 4717
rect 2889 4691 2915 4717
rect 2915 4691 2916 4717
rect 2888 4690 2916 4691
rect 2940 4717 2968 4718
rect 2940 4691 2941 4717
rect 2941 4691 2967 4717
rect 2967 4691 2968 4717
rect 2940 4690 2968 4691
rect 2992 4717 3020 4718
rect 2992 4691 2993 4717
rect 2993 4691 3019 4717
rect 3019 4691 3020 4717
rect 2992 4690 3020 4691
rect 3044 4717 3072 4718
rect 3044 4691 3045 4717
rect 3045 4691 3071 4717
rect 3071 4691 3072 4717
rect 3044 4690 3072 4691
rect 3096 4717 3124 4718
rect 3096 4691 3097 4717
rect 3097 4691 3123 4717
rect 3123 4691 3124 4717
rect 3096 4690 3124 4691
rect 3148 4717 3176 4718
rect 3148 4691 3149 4717
rect 3149 4691 3175 4717
rect 3175 4691 3176 4717
rect 3148 4690 3176 4691
rect 1078 4521 1106 4522
rect 1078 4495 1079 4521
rect 1079 4495 1105 4521
rect 1105 4495 1106 4521
rect 1078 4494 1106 4495
rect 1358 4521 1386 4522
rect 1358 4495 1359 4521
rect 1359 4495 1385 4521
rect 1385 4495 1386 4521
rect 1358 4494 1386 4495
rect 1028 4325 1056 4326
rect 1028 4299 1029 4325
rect 1029 4299 1055 4325
rect 1055 4299 1056 4325
rect 1028 4298 1056 4299
rect 1080 4325 1108 4326
rect 1080 4299 1081 4325
rect 1081 4299 1107 4325
rect 1107 4299 1108 4325
rect 1080 4298 1108 4299
rect 1132 4325 1160 4326
rect 1132 4299 1133 4325
rect 1133 4299 1159 4325
rect 1159 4299 1160 4325
rect 1132 4298 1160 4299
rect 1184 4325 1212 4326
rect 1184 4299 1185 4325
rect 1185 4299 1211 4325
rect 1211 4299 1212 4325
rect 1184 4298 1212 4299
rect 1236 4325 1264 4326
rect 1236 4299 1237 4325
rect 1237 4299 1263 4325
rect 1263 4299 1264 4325
rect 1236 4298 1264 4299
rect 1288 4325 1316 4326
rect 1288 4299 1289 4325
rect 1289 4299 1315 4325
rect 1315 4299 1316 4325
rect 1288 4298 1316 4299
rect 910 4158 938 4186
rect 2888 3933 2916 3934
rect 2888 3907 2889 3933
rect 2889 3907 2915 3933
rect 2915 3907 2916 3933
rect 2888 3906 2916 3907
rect 2940 3933 2968 3934
rect 2940 3907 2941 3933
rect 2941 3907 2967 3933
rect 2967 3907 2968 3933
rect 2940 3906 2968 3907
rect 2992 3933 3020 3934
rect 2992 3907 2993 3933
rect 2993 3907 3019 3933
rect 3019 3907 3020 3933
rect 2992 3906 3020 3907
rect 3044 3933 3072 3934
rect 3044 3907 3045 3933
rect 3045 3907 3071 3933
rect 3071 3907 3072 3933
rect 3044 3906 3072 3907
rect 3096 3933 3124 3934
rect 3096 3907 3097 3933
rect 3097 3907 3123 3933
rect 3123 3907 3124 3933
rect 3096 3906 3124 3907
rect 3148 3933 3176 3934
rect 3148 3907 3149 3933
rect 3149 3907 3175 3933
rect 3175 3907 3176 3933
rect 3148 3906 3176 3907
rect 1028 3541 1056 3542
rect 1028 3515 1029 3541
rect 1029 3515 1055 3541
rect 1055 3515 1056 3541
rect 1028 3514 1056 3515
rect 1080 3541 1108 3542
rect 1080 3515 1081 3541
rect 1081 3515 1107 3541
rect 1107 3515 1108 3541
rect 1080 3514 1108 3515
rect 1132 3541 1160 3542
rect 1132 3515 1133 3541
rect 1133 3515 1159 3541
rect 1159 3515 1160 3541
rect 1132 3514 1160 3515
rect 1184 3541 1212 3542
rect 1184 3515 1185 3541
rect 1185 3515 1211 3541
rect 1211 3515 1212 3541
rect 1184 3514 1212 3515
rect 1236 3541 1264 3542
rect 1236 3515 1237 3541
rect 1237 3515 1263 3541
rect 1263 3515 1264 3541
rect 1236 3514 1264 3515
rect 1288 3541 1316 3542
rect 1288 3515 1289 3541
rect 1289 3515 1315 3541
rect 1315 3515 1316 3541
rect 1288 3514 1316 3515
rect 2888 3149 2916 3150
rect 2888 3123 2889 3149
rect 2889 3123 2915 3149
rect 2915 3123 2916 3149
rect 2888 3122 2916 3123
rect 2940 3149 2968 3150
rect 2940 3123 2941 3149
rect 2941 3123 2967 3149
rect 2967 3123 2968 3149
rect 2940 3122 2968 3123
rect 2992 3149 3020 3150
rect 2992 3123 2993 3149
rect 2993 3123 3019 3149
rect 3019 3123 3020 3149
rect 2992 3122 3020 3123
rect 3044 3149 3072 3150
rect 3044 3123 3045 3149
rect 3045 3123 3071 3149
rect 3071 3123 3072 3149
rect 3044 3122 3072 3123
rect 3096 3149 3124 3150
rect 3096 3123 3097 3149
rect 3097 3123 3123 3149
rect 3123 3123 3124 3149
rect 3096 3122 3124 3123
rect 3148 3149 3176 3150
rect 3148 3123 3149 3149
rect 3149 3123 3175 3149
rect 3175 3123 3176 3149
rect 3148 3122 3176 3123
rect 1028 2757 1056 2758
rect 1028 2731 1029 2757
rect 1029 2731 1055 2757
rect 1055 2731 1056 2757
rect 1028 2730 1056 2731
rect 1080 2757 1108 2758
rect 1080 2731 1081 2757
rect 1081 2731 1107 2757
rect 1107 2731 1108 2757
rect 1080 2730 1108 2731
rect 1132 2757 1160 2758
rect 1132 2731 1133 2757
rect 1133 2731 1159 2757
rect 1159 2731 1160 2757
rect 1132 2730 1160 2731
rect 1184 2757 1212 2758
rect 1184 2731 1185 2757
rect 1185 2731 1211 2757
rect 1211 2731 1212 2757
rect 1184 2730 1212 2731
rect 1236 2757 1264 2758
rect 1236 2731 1237 2757
rect 1237 2731 1263 2757
rect 1263 2731 1264 2757
rect 1236 2730 1264 2731
rect 1288 2757 1316 2758
rect 1288 2731 1289 2757
rect 1289 2731 1315 2757
rect 1315 2731 1316 2757
rect 1288 2730 1316 2731
rect 2888 2365 2916 2366
rect 2888 2339 2889 2365
rect 2889 2339 2915 2365
rect 2915 2339 2916 2365
rect 2888 2338 2916 2339
rect 2940 2365 2968 2366
rect 2940 2339 2941 2365
rect 2941 2339 2967 2365
rect 2967 2339 2968 2365
rect 2940 2338 2968 2339
rect 2992 2365 3020 2366
rect 2992 2339 2993 2365
rect 2993 2339 3019 2365
rect 3019 2339 3020 2365
rect 2992 2338 3020 2339
rect 3044 2365 3072 2366
rect 3044 2339 3045 2365
rect 3045 2339 3071 2365
rect 3071 2339 3072 2365
rect 3044 2338 3072 2339
rect 3096 2365 3124 2366
rect 3096 2339 3097 2365
rect 3097 2339 3123 2365
rect 3123 2339 3124 2365
rect 3096 2338 3124 2339
rect 3148 2365 3176 2366
rect 3148 2339 3149 2365
rect 3149 2339 3175 2365
rect 3175 2339 3176 2365
rect 3148 2338 3176 2339
rect 1028 1973 1056 1974
rect 1028 1947 1029 1973
rect 1029 1947 1055 1973
rect 1055 1947 1056 1973
rect 1028 1946 1056 1947
rect 1080 1973 1108 1974
rect 1080 1947 1081 1973
rect 1081 1947 1107 1973
rect 1107 1947 1108 1973
rect 1080 1946 1108 1947
rect 1132 1973 1160 1974
rect 1132 1947 1133 1973
rect 1133 1947 1159 1973
rect 1159 1947 1160 1973
rect 1132 1946 1160 1947
rect 1184 1973 1212 1974
rect 1184 1947 1185 1973
rect 1185 1947 1211 1973
rect 1211 1947 1212 1973
rect 1184 1946 1212 1947
rect 1236 1973 1264 1974
rect 1236 1947 1237 1973
rect 1237 1947 1263 1973
rect 1263 1947 1264 1973
rect 1236 1946 1264 1947
rect 1288 1973 1316 1974
rect 1288 1947 1289 1973
rect 1289 1947 1315 1973
rect 1315 1947 1316 1973
rect 1288 1946 1316 1947
rect 2888 1581 2916 1582
rect 2888 1555 2889 1581
rect 2889 1555 2915 1581
rect 2915 1555 2916 1581
rect 2888 1554 2916 1555
rect 2940 1581 2968 1582
rect 2940 1555 2941 1581
rect 2941 1555 2967 1581
rect 2967 1555 2968 1581
rect 2940 1554 2968 1555
rect 2992 1581 3020 1582
rect 2992 1555 2993 1581
rect 2993 1555 3019 1581
rect 3019 1555 3020 1581
rect 2992 1554 3020 1555
rect 3044 1581 3072 1582
rect 3044 1555 3045 1581
rect 3045 1555 3071 1581
rect 3071 1555 3072 1581
rect 3044 1554 3072 1555
rect 3096 1581 3124 1582
rect 3096 1555 3097 1581
rect 3097 1555 3123 1581
rect 3123 1555 3124 1581
rect 3096 1554 3124 1555
rect 3148 1581 3176 1582
rect 3148 1555 3149 1581
rect 3149 1555 3175 1581
rect 3175 1555 3176 1581
rect 3148 1554 3176 1555
rect 10878 4886 10906 4914
rect 12502 5249 12530 5250
rect 12502 5223 12503 5249
rect 12503 5223 12529 5249
rect 12529 5223 12530 5249
rect 12502 5222 12530 5223
rect 12838 5222 12866 5250
rect 12446 5166 12474 5194
rect 11886 4913 11914 4914
rect 11886 4887 11887 4913
rect 11887 4887 11913 4913
rect 11913 4887 11914 4913
rect 11886 4886 11914 4887
rect 12278 4774 12306 4802
rect 11718 4494 11746 4522
rect 16030 6089 16058 6090
rect 16030 6063 16031 6089
rect 16031 6063 16057 6089
rect 16057 6063 16058 6089
rect 16030 6062 16058 6063
rect 16254 6089 16282 6090
rect 16254 6063 16255 6089
rect 16255 6063 16281 6089
rect 16281 6063 16282 6089
rect 16254 6062 16282 6063
rect 19028 5893 19056 5894
rect 19028 5867 19029 5893
rect 19029 5867 19055 5893
rect 19055 5867 19056 5893
rect 19028 5866 19056 5867
rect 19080 5893 19108 5894
rect 19080 5867 19081 5893
rect 19081 5867 19107 5893
rect 19107 5867 19108 5893
rect 19080 5866 19108 5867
rect 19132 5893 19160 5894
rect 19132 5867 19133 5893
rect 19133 5867 19159 5893
rect 19159 5867 19160 5893
rect 19132 5866 19160 5867
rect 19184 5893 19212 5894
rect 19184 5867 19185 5893
rect 19185 5867 19211 5893
rect 19211 5867 19212 5893
rect 19184 5866 19212 5867
rect 19236 5893 19264 5894
rect 19236 5867 19237 5893
rect 19237 5867 19263 5893
rect 19263 5867 19264 5893
rect 19236 5866 19264 5867
rect 19288 5893 19316 5894
rect 19288 5867 19289 5893
rect 19289 5867 19315 5893
rect 19315 5867 19316 5893
rect 19288 5866 19316 5867
rect 22246 5558 22274 5586
rect 20888 5501 20916 5502
rect 20888 5475 20889 5501
rect 20889 5475 20915 5501
rect 20915 5475 20916 5501
rect 20888 5474 20916 5475
rect 20940 5501 20968 5502
rect 20940 5475 20941 5501
rect 20941 5475 20967 5501
rect 20967 5475 20968 5501
rect 20940 5474 20968 5475
rect 20992 5501 21020 5502
rect 20992 5475 20993 5501
rect 20993 5475 21019 5501
rect 21019 5475 21020 5501
rect 20992 5474 21020 5475
rect 21044 5501 21072 5502
rect 21044 5475 21045 5501
rect 21045 5475 21071 5501
rect 21071 5475 21072 5501
rect 21044 5474 21072 5475
rect 21096 5501 21124 5502
rect 21096 5475 21097 5501
rect 21097 5475 21123 5501
rect 21123 5475 21124 5501
rect 21096 5474 21124 5475
rect 21148 5501 21176 5502
rect 21148 5475 21149 5501
rect 21149 5475 21175 5501
rect 21175 5475 21176 5501
rect 21148 5474 21176 5475
rect 14294 5166 14322 5194
rect 19028 5109 19056 5110
rect 19028 5083 19029 5109
rect 19029 5083 19055 5109
rect 19055 5083 19056 5109
rect 19028 5082 19056 5083
rect 19080 5109 19108 5110
rect 19080 5083 19081 5109
rect 19081 5083 19107 5109
rect 19107 5083 19108 5109
rect 19080 5082 19108 5083
rect 19132 5109 19160 5110
rect 19132 5083 19133 5109
rect 19133 5083 19159 5109
rect 19159 5083 19160 5109
rect 19132 5082 19160 5083
rect 19184 5109 19212 5110
rect 19184 5083 19185 5109
rect 19185 5083 19211 5109
rect 19211 5083 19212 5109
rect 19184 5082 19212 5083
rect 19236 5109 19264 5110
rect 19236 5083 19237 5109
rect 19237 5083 19263 5109
rect 19263 5083 19264 5109
rect 19236 5082 19264 5083
rect 19288 5109 19316 5110
rect 19288 5083 19289 5109
rect 19289 5083 19315 5109
rect 19315 5083 19316 5109
rect 19288 5082 19316 5083
rect 13566 4801 13594 4802
rect 13566 4775 13567 4801
rect 13567 4775 13593 4801
rect 13593 4775 13594 4801
rect 13566 4774 13594 4775
rect 18830 4774 18858 4802
rect 18662 1694 18690 1722
rect 20888 4717 20916 4718
rect 20888 4691 20889 4717
rect 20889 4691 20915 4717
rect 20915 4691 20916 4717
rect 20888 4690 20916 4691
rect 20940 4717 20968 4718
rect 20940 4691 20941 4717
rect 20941 4691 20967 4717
rect 20967 4691 20968 4717
rect 20940 4690 20968 4691
rect 20992 4717 21020 4718
rect 20992 4691 20993 4717
rect 20993 4691 21019 4717
rect 21019 4691 21020 4717
rect 20992 4690 21020 4691
rect 21044 4717 21072 4718
rect 21044 4691 21045 4717
rect 21045 4691 21071 4717
rect 21071 4691 21072 4717
rect 21044 4690 21072 4691
rect 21096 4717 21124 4718
rect 21096 4691 21097 4717
rect 21097 4691 21123 4717
rect 21123 4691 21124 4717
rect 21096 4690 21124 4691
rect 21148 4717 21176 4718
rect 21148 4691 21149 4717
rect 21149 4691 21175 4717
rect 21175 4691 21176 4717
rect 21148 4690 21176 4691
rect 19028 4325 19056 4326
rect 19028 4299 19029 4325
rect 19029 4299 19055 4325
rect 19055 4299 19056 4325
rect 19028 4298 19056 4299
rect 19080 4325 19108 4326
rect 19080 4299 19081 4325
rect 19081 4299 19107 4325
rect 19107 4299 19108 4325
rect 19080 4298 19108 4299
rect 19132 4325 19160 4326
rect 19132 4299 19133 4325
rect 19133 4299 19159 4325
rect 19159 4299 19160 4325
rect 19132 4298 19160 4299
rect 19184 4325 19212 4326
rect 19184 4299 19185 4325
rect 19185 4299 19211 4325
rect 19211 4299 19212 4325
rect 19184 4298 19212 4299
rect 19236 4325 19264 4326
rect 19236 4299 19237 4325
rect 19237 4299 19263 4325
rect 19263 4299 19264 4325
rect 19236 4298 19264 4299
rect 19288 4325 19316 4326
rect 19288 4299 19289 4325
rect 19289 4299 19315 4325
rect 19315 4299 19316 4325
rect 19288 4298 19316 4299
rect 20888 3933 20916 3934
rect 20888 3907 20889 3933
rect 20889 3907 20915 3933
rect 20915 3907 20916 3933
rect 20888 3906 20916 3907
rect 20940 3933 20968 3934
rect 20940 3907 20941 3933
rect 20941 3907 20967 3933
rect 20967 3907 20968 3933
rect 20940 3906 20968 3907
rect 20992 3933 21020 3934
rect 20992 3907 20993 3933
rect 20993 3907 21019 3933
rect 21019 3907 21020 3933
rect 20992 3906 21020 3907
rect 21044 3933 21072 3934
rect 21044 3907 21045 3933
rect 21045 3907 21071 3933
rect 21071 3907 21072 3933
rect 21044 3906 21072 3907
rect 21096 3933 21124 3934
rect 21096 3907 21097 3933
rect 21097 3907 21123 3933
rect 21123 3907 21124 3933
rect 21096 3906 21124 3907
rect 21148 3933 21176 3934
rect 21148 3907 21149 3933
rect 21149 3907 21175 3933
rect 21175 3907 21176 3933
rect 21148 3906 21176 3907
rect 19028 3541 19056 3542
rect 19028 3515 19029 3541
rect 19029 3515 19055 3541
rect 19055 3515 19056 3541
rect 19028 3514 19056 3515
rect 19080 3541 19108 3542
rect 19080 3515 19081 3541
rect 19081 3515 19107 3541
rect 19107 3515 19108 3541
rect 19080 3514 19108 3515
rect 19132 3541 19160 3542
rect 19132 3515 19133 3541
rect 19133 3515 19159 3541
rect 19159 3515 19160 3541
rect 19132 3514 19160 3515
rect 19184 3541 19212 3542
rect 19184 3515 19185 3541
rect 19185 3515 19211 3541
rect 19211 3515 19212 3541
rect 19184 3514 19212 3515
rect 19236 3541 19264 3542
rect 19236 3515 19237 3541
rect 19237 3515 19263 3541
rect 19263 3515 19264 3541
rect 19236 3514 19264 3515
rect 19288 3541 19316 3542
rect 19288 3515 19289 3541
rect 19289 3515 19315 3541
rect 19315 3515 19316 3541
rect 19288 3514 19316 3515
rect 20888 3149 20916 3150
rect 20888 3123 20889 3149
rect 20889 3123 20915 3149
rect 20915 3123 20916 3149
rect 20888 3122 20916 3123
rect 20940 3149 20968 3150
rect 20940 3123 20941 3149
rect 20941 3123 20967 3149
rect 20967 3123 20968 3149
rect 20940 3122 20968 3123
rect 20992 3149 21020 3150
rect 20992 3123 20993 3149
rect 20993 3123 21019 3149
rect 21019 3123 21020 3149
rect 20992 3122 21020 3123
rect 21044 3149 21072 3150
rect 21044 3123 21045 3149
rect 21045 3123 21071 3149
rect 21071 3123 21072 3149
rect 21044 3122 21072 3123
rect 21096 3149 21124 3150
rect 21096 3123 21097 3149
rect 21097 3123 21123 3149
rect 21123 3123 21124 3149
rect 21096 3122 21124 3123
rect 21148 3149 21176 3150
rect 21148 3123 21149 3149
rect 21149 3123 21175 3149
rect 21175 3123 21176 3149
rect 21148 3122 21176 3123
rect 19028 2757 19056 2758
rect 19028 2731 19029 2757
rect 19029 2731 19055 2757
rect 19055 2731 19056 2757
rect 19028 2730 19056 2731
rect 19080 2757 19108 2758
rect 19080 2731 19081 2757
rect 19081 2731 19107 2757
rect 19107 2731 19108 2757
rect 19080 2730 19108 2731
rect 19132 2757 19160 2758
rect 19132 2731 19133 2757
rect 19133 2731 19159 2757
rect 19159 2731 19160 2757
rect 19132 2730 19160 2731
rect 19184 2757 19212 2758
rect 19184 2731 19185 2757
rect 19185 2731 19211 2757
rect 19211 2731 19212 2757
rect 19184 2730 19212 2731
rect 19236 2757 19264 2758
rect 19236 2731 19237 2757
rect 19237 2731 19263 2757
rect 19263 2731 19264 2757
rect 19236 2730 19264 2731
rect 19288 2757 19316 2758
rect 19288 2731 19289 2757
rect 19289 2731 19315 2757
rect 19315 2731 19316 2757
rect 19288 2730 19316 2731
rect 20888 2365 20916 2366
rect 20888 2339 20889 2365
rect 20889 2339 20915 2365
rect 20915 2339 20916 2365
rect 20888 2338 20916 2339
rect 20940 2365 20968 2366
rect 20940 2339 20941 2365
rect 20941 2339 20967 2365
rect 20967 2339 20968 2365
rect 20940 2338 20968 2339
rect 20992 2365 21020 2366
rect 20992 2339 20993 2365
rect 20993 2339 21019 2365
rect 21019 2339 21020 2365
rect 20992 2338 21020 2339
rect 21044 2365 21072 2366
rect 21044 2339 21045 2365
rect 21045 2339 21071 2365
rect 21071 2339 21072 2365
rect 21044 2338 21072 2339
rect 21096 2365 21124 2366
rect 21096 2339 21097 2365
rect 21097 2339 21123 2365
rect 21123 2339 21124 2365
rect 21096 2338 21124 2339
rect 21148 2365 21176 2366
rect 21148 2339 21149 2365
rect 21149 2339 21175 2365
rect 21175 2339 21176 2365
rect 21148 2338 21176 2339
rect 19028 1973 19056 1974
rect 19028 1947 19029 1973
rect 19029 1947 19055 1973
rect 19055 1947 19056 1973
rect 19028 1946 19056 1947
rect 19080 1973 19108 1974
rect 19080 1947 19081 1973
rect 19081 1947 19107 1973
rect 19107 1947 19108 1973
rect 19080 1946 19108 1947
rect 19132 1973 19160 1974
rect 19132 1947 19133 1973
rect 19133 1947 19159 1973
rect 19159 1947 19160 1973
rect 19132 1946 19160 1947
rect 19184 1973 19212 1974
rect 19184 1947 19185 1973
rect 19185 1947 19211 1973
rect 19211 1947 19212 1973
rect 19184 1946 19212 1947
rect 19236 1973 19264 1974
rect 19236 1947 19237 1973
rect 19237 1947 19263 1973
rect 19263 1947 19264 1973
rect 19236 1946 19264 1947
rect 19288 1973 19316 1974
rect 19288 1947 19289 1973
rect 19289 1947 19315 1973
rect 19315 1947 19316 1973
rect 19288 1946 19316 1947
rect 18998 1721 19026 1722
rect 18998 1695 18999 1721
rect 18999 1695 19025 1721
rect 19025 1695 19026 1721
rect 18998 1694 19026 1695
rect 20888 1581 20916 1582
rect 20888 1555 20889 1581
rect 20889 1555 20915 1581
rect 20915 1555 20916 1581
rect 20888 1554 20916 1555
rect 20940 1581 20968 1582
rect 20940 1555 20941 1581
rect 20941 1555 20967 1581
rect 20967 1555 20968 1581
rect 20940 1554 20968 1555
rect 20992 1581 21020 1582
rect 20992 1555 20993 1581
rect 20993 1555 21019 1581
rect 21019 1555 21020 1581
rect 20992 1554 21020 1555
rect 21044 1581 21072 1582
rect 21044 1555 21045 1581
rect 21045 1555 21071 1581
rect 21071 1555 21072 1581
rect 21044 1554 21072 1555
rect 21096 1581 21124 1582
rect 21096 1555 21097 1581
rect 21097 1555 21123 1581
rect 21123 1555 21124 1581
rect 21096 1554 21124 1555
rect 21148 1581 21176 1582
rect 21148 1555 21149 1581
rect 21149 1555 21175 1581
rect 21175 1555 21176 1581
rect 21148 1554 21176 1555
<< metal3 >>
rect 1023 23114 1028 23142
rect 1056 23114 1080 23142
rect 1108 23114 1132 23142
rect 1160 23114 1184 23142
rect 1212 23114 1236 23142
rect 1264 23114 1288 23142
rect 1316 23114 1321 23142
rect 19023 23114 19028 23142
rect 19056 23114 19080 23142
rect 19108 23114 19132 23142
rect 19160 23114 19184 23142
rect 19212 23114 19236 23142
rect 19264 23114 19288 23142
rect 19316 23114 19321 23142
rect 2883 22722 2888 22750
rect 2916 22722 2940 22750
rect 2968 22722 2992 22750
rect 3020 22722 3044 22750
rect 3072 22722 3096 22750
rect 3124 22722 3148 22750
rect 3176 22722 3181 22750
rect 20883 22722 20888 22750
rect 20916 22722 20940 22750
rect 20968 22722 20992 22750
rect 21020 22722 21044 22750
rect 21072 22722 21096 22750
rect 21124 22722 21148 22750
rect 21176 22722 21181 22750
rect 1023 22330 1028 22358
rect 1056 22330 1080 22358
rect 1108 22330 1132 22358
rect 1160 22330 1184 22358
rect 1212 22330 1236 22358
rect 1264 22330 1288 22358
rect 1316 22330 1321 22358
rect 19023 22330 19028 22358
rect 19056 22330 19080 22358
rect 19108 22330 19132 22358
rect 19160 22330 19184 22358
rect 19212 22330 19236 22358
rect 19264 22330 19288 22358
rect 19316 22330 19321 22358
rect 2883 21938 2888 21966
rect 2916 21938 2940 21966
rect 2968 21938 2992 21966
rect 3020 21938 3044 21966
rect 3072 21938 3096 21966
rect 3124 21938 3148 21966
rect 3176 21938 3181 21966
rect 20883 21938 20888 21966
rect 20916 21938 20940 21966
rect 20968 21938 20992 21966
rect 21020 21938 21044 21966
rect 21072 21938 21096 21966
rect 21124 21938 21148 21966
rect 21176 21938 21181 21966
rect 1023 21546 1028 21574
rect 1056 21546 1080 21574
rect 1108 21546 1132 21574
rect 1160 21546 1184 21574
rect 1212 21546 1236 21574
rect 1264 21546 1288 21574
rect 1316 21546 1321 21574
rect 19023 21546 19028 21574
rect 19056 21546 19080 21574
rect 19108 21546 19132 21574
rect 19160 21546 19184 21574
rect 19212 21546 19236 21574
rect 19264 21546 19288 21574
rect 19316 21546 19321 21574
rect 2883 21154 2888 21182
rect 2916 21154 2940 21182
rect 2968 21154 2992 21182
rect 3020 21154 3044 21182
rect 3072 21154 3096 21182
rect 3124 21154 3148 21182
rect 3176 21154 3181 21182
rect 20883 21154 20888 21182
rect 20916 21154 20940 21182
rect 20968 21154 20992 21182
rect 21020 21154 21044 21182
rect 21072 21154 21096 21182
rect 21124 21154 21148 21182
rect 21176 21154 21181 21182
rect 196 20804 910 20818
rect -480 20790 910 20804
rect 938 20790 943 20818
rect -480 20692 240 20790
rect 1023 20762 1028 20790
rect 1056 20762 1080 20790
rect 1108 20762 1132 20790
rect 1160 20762 1184 20790
rect 1212 20762 1236 20790
rect 1264 20762 1288 20790
rect 1316 20762 1321 20790
rect 19023 20762 19028 20790
rect 19056 20762 19080 20790
rect 19108 20762 19132 20790
rect 19160 20762 19184 20790
rect 19212 20762 19236 20790
rect 19264 20762 19288 20790
rect 19316 20762 19321 20790
rect 2883 20370 2888 20398
rect 2916 20370 2940 20398
rect 2968 20370 2992 20398
rect 3020 20370 3044 20398
rect 3072 20370 3096 20398
rect 3124 20370 3148 20398
rect 3176 20370 3181 20398
rect 20883 20370 20888 20398
rect 20916 20370 20940 20398
rect 20968 20370 20992 20398
rect 21020 20370 21044 20398
rect 21072 20370 21096 20398
rect 21124 20370 21148 20398
rect 21176 20370 21181 20398
rect 1023 19978 1028 20006
rect 1056 19978 1080 20006
rect 1108 19978 1132 20006
rect 1160 19978 1184 20006
rect 1212 19978 1236 20006
rect 1264 19978 1288 20006
rect 1316 19978 1321 20006
rect 19023 19978 19028 20006
rect 19056 19978 19080 20006
rect 19108 19978 19132 20006
rect 19160 19978 19184 20006
rect 19212 19978 19236 20006
rect 19264 19978 19288 20006
rect 19316 19978 19321 20006
rect 2883 19586 2888 19614
rect 2916 19586 2940 19614
rect 2968 19586 2992 19614
rect 3020 19586 3044 19614
rect 3072 19586 3096 19614
rect 3124 19586 3148 19614
rect 3176 19586 3181 19614
rect 20883 19586 20888 19614
rect 20916 19586 20940 19614
rect 20968 19586 20992 19614
rect 21020 19586 21044 19614
rect 21072 19586 21096 19614
rect 21124 19586 21148 19614
rect 21176 19586 21181 19614
rect 1023 19194 1028 19222
rect 1056 19194 1080 19222
rect 1108 19194 1132 19222
rect 1160 19194 1184 19222
rect 1212 19194 1236 19222
rect 1264 19194 1288 19222
rect 1316 19194 1321 19222
rect 19023 19194 19028 19222
rect 19056 19194 19080 19222
rect 19108 19194 19132 19222
rect 19160 19194 19184 19222
rect 19212 19194 19236 19222
rect 19264 19194 19288 19222
rect 19316 19194 19321 19222
rect 2883 18802 2888 18830
rect 2916 18802 2940 18830
rect 2968 18802 2992 18830
rect 3020 18802 3044 18830
rect 3072 18802 3096 18830
rect 3124 18802 3148 18830
rect 3176 18802 3181 18830
rect 20883 18802 20888 18830
rect 20916 18802 20940 18830
rect 20968 18802 20992 18830
rect 21020 18802 21044 18830
rect 21072 18802 21096 18830
rect 21124 18802 21148 18830
rect 21176 18802 21181 18830
rect 1023 18410 1028 18438
rect 1056 18410 1080 18438
rect 1108 18410 1132 18438
rect 1160 18410 1184 18438
rect 1212 18410 1236 18438
rect 1264 18410 1288 18438
rect 1316 18410 1321 18438
rect 19023 18410 19028 18438
rect 19056 18410 19080 18438
rect 19108 18410 19132 18438
rect 19160 18410 19184 18438
rect 19212 18410 19236 18438
rect 19264 18410 19288 18438
rect 19316 18410 19321 18438
rect 2883 18018 2888 18046
rect 2916 18018 2940 18046
rect 2968 18018 2992 18046
rect 3020 18018 3044 18046
rect 3072 18018 3096 18046
rect 3124 18018 3148 18046
rect 3176 18018 3181 18046
rect 20883 18018 20888 18046
rect 20916 18018 20940 18046
rect 20968 18018 20992 18046
rect 21020 18018 21044 18046
rect 21072 18018 21096 18046
rect 21124 18018 21148 18046
rect 21176 18018 21181 18046
rect 1023 17626 1028 17654
rect 1056 17626 1080 17654
rect 1108 17626 1132 17654
rect 1160 17626 1184 17654
rect 1212 17626 1236 17654
rect 1264 17626 1288 17654
rect 1316 17626 1321 17654
rect 19023 17626 19028 17654
rect 19056 17626 19080 17654
rect 19108 17626 19132 17654
rect 19160 17626 19184 17654
rect 19212 17626 19236 17654
rect 19264 17626 19288 17654
rect 19316 17626 19321 17654
rect 2883 17234 2888 17262
rect 2916 17234 2940 17262
rect 2968 17234 2992 17262
rect 3020 17234 3044 17262
rect 3072 17234 3096 17262
rect 3124 17234 3148 17262
rect 3176 17234 3181 17262
rect 20883 17234 20888 17262
rect 20916 17234 20940 17262
rect 20968 17234 20992 17262
rect 21020 17234 21044 17262
rect 21072 17234 21096 17262
rect 21124 17234 21148 17262
rect 21176 17234 21181 17262
rect 1023 16842 1028 16870
rect 1056 16842 1080 16870
rect 1108 16842 1132 16870
rect 1160 16842 1184 16870
rect 1212 16842 1236 16870
rect 1264 16842 1288 16870
rect 1316 16842 1321 16870
rect 19023 16842 19028 16870
rect 19056 16842 19080 16870
rect 19108 16842 19132 16870
rect 19160 16842 19184 16870
rect 19212 16842 19236 16870
rect 19264 16842 19288 16870
rect 19316 16842 19321 16870
rect 2883 16450 2888 16478
rect 2916 16450 2940 16478
rect 2968 16450 2992 16478
rect 3020 16450 3044 16478
rect 3072 16450 3096 16478
rect 3124 16450 3148 16478
rect 3176 16450 3181 16478
rect 20883 16450 20888 16478
rect 20916 16450 20940 16478
rect 20968 16450 20992 16478
rect 21020 16450 21044 16478
rect 21072 16450 21096 16478
rect 21124 16450 21148 16478
rect 21176 16450 21181 16478
rect 1023 16058 1028 16086
rect 1056 16058 1080 16086
rect 1108 16058 1132 16086
rect 1160 16058 1184 16086
rect 1212 16058 1236 16086
rect 1264 16058 1288 16086
rect 1316 16058 1321 16086
rect 19023 16058 19028 16086
rect 19056 16058 19080 16086
rect 19108 16058 19132 16086
rect 19160 16058 19184 16086
rect 19212 16058 19236 16086
rect 19264 16058 19288 16086
rect 19316 16058 19321 16086
rect 2883 15666 2888 15694
rect 2916 15666 2940 15694
rect 2968 15666 2992 15694
rect 3020 15666 3044 15694
rect 3072 15666 3096 15694
rect 3124 15666 3148 15694
rect 3176 15666 3181 15694
rect 20883 15666 20888 15694
rect 20916 15666 20940 15694
rect 20968 15666 20992 15694
rect 21020 15666 21044 15694
rect 21072 15666 21096 15694
rect 21124 15666 21148 15694
rect 21176 15666 21181 15694
rect 1023 15274 1028 15302
rect 1056 15274 1080 15302
rect 1108 15274 1132 15302
rect 1160 15274 1184 15302
rect 1212 15274 1236 15302
rect 1264 15274 1288 15302
rect 1316 15274 1321 15302
rect 19023 15274 19028 15302
rect 19056 15274 19080 15302
rect 19108 15274 19132 15302
rect 19160 15274 19184 15302
rect 19212 15274 19236 15302
rect 19264 15274 19288 15302
rect 19316 15274 19321 15302
rect 2883 14882 2888 14910
rect 2916 14882 2940 14910
rect 2968 14882 2992 14910
rect 3020 14882 3044 14910
rect 3072 14882 3096 14910
rect 3124 14882 3148 14910
rect 3176 14882 3181 14910
rect 20883 14882 20888 14910
rect 20916 14882 20940 14910
rect 20968 14882 20992 14910
rect 21020 14882 21044 14910
rect 21072 14882 21096 14910
rect 21124 14882 21148 14910
rect 21176 14882 21181 14910
rect 1023 14490 1028 14518
rect 1056 14490 1080 14518
rect 1108 14490 1132 14518
rect 1160 14490 1184 14518
rect 1212 14490 1236 14518
rect 1264 14490 1288 14518
rect 1316 14490 1321 14518
rect 19023 14490 19028 14518
rect 19056 14490 19080 14518
rect 19108 14490 19132 14518
rect 19160 14490 19184 14518
rect 19212 14490 19236 14518
rect 19264 14490 19288 14518
rect 19316 14490 19321 14518
rect 2883 14098 2888 14126
rect 2916 14098 2940 14126
rect 2968 14098 2992 14126
rect 3020 14098 3044 14126
rect 3072 14098 3096 14126
rect 3124 14098 3148 14126
rect 3176 14098 3181 14126
rect 20883 14098 20888 14126
rect 20916 14098 20940 14126
rect 20968 14098 20992 14126
rect 21020 14098 21044 14126
rect 21072 14098 21096 14126
rect 21124 14098 21148 14126
rect 21176 14098 21181 14126
rect 1023 13706 1028 13734
rect 1056 13706 1080 13734
rect 1108 13706 1132 13734
rect 1160 13706 1184 13734
rect 1212 13706 1236 13734
rect 1264 13706 1288 13734
rect 1316 13706 1321 13734
rect 19023 13706 19028 13734
rect 19056 13706 19080 13734
rect 19108 13706 19132 13734
rect 19160 13706 19184 13734
rect 19212 13706 19236 13734
rect 19264 13706 19288 13734
rect 19316 13706 19321 13734
rect 2883 13314 2888 13342
rect 2916 13314 2940 13342
rect 2968 13314 2992 13342
rect 3020 13314 3044 13342
rect 3072 13314 3096 13342
rect 3124 13314 3148 13342
rect 3176 13314 3181 13342
rect 20883 13314 20888 13342
rect 20916 13314 20940 13342
rect 20968 13314 20992 13342
rect 21020 13314 21044 13342
rect 21072 13314 21096 13342
rect 21124 13314 21148 13342
rect 21176 13314 21181 13342
rect 1023 12922 1028 12950
rect 1056 12922 1080 12950
rect 1108 12922 1132 12950
rect 1160 12922 1184 12950
rect 1212 12922 1236 12950
rect 1264 12922 1288 12950
rect 1316 12922 1321 12950
rect 19023 12922 19028 12950
rect 19056 12922 19080 12950
rect 19108 12922 19132 12950
rect 19160 12922 19184 12950
rect 19212 12922 19236 12950
rect 19264 12922 19288 12950
rect 19316 12922 19321 12950
rect 2883 12530 2888 12558
rect 2916 12530 2940 12558
rect 2968 12530 2992 12558
rect 3020 12530 3044 12558
rect 3072 12530 3096 12558
rect 3124 12530 3148 12558
rect 3176 12530 3181 12558
rect 20883 12530 20888 12558
rect 20916 12530 20940 12558
rect 20968 12530 20992 12558
rect 21020 12530 21044 12558
rect 21072 12530 21096 12558
rect 21124 12530 21148 12558
rect 21176 12530 21181 12558
rect 196 12516 910 12530
rect -480 12502 910 12516
rect 938 12502 943 12530
rect -480 12404 240 12502
rect 24760 12474 25480 12516
rect 22241 12446 22246 12474
rect 22274 12446 25480 12474
rect 24760 12404 25480 12446
rect 1023 12138 1028 12166
rect 1056 12138 1080 12166
rect 1108 12138 1132 12166
rect 1160 12138 1184 12166
rect 1212 12138 1236 12166
rect 1264 12138 1288 12166
rect 1316 12138 1321 12166
rect 19023 12138 19028 12166
rect 19056 12138 19080 12166
rect 19108 12138 19132 12166
rect 19160 12138 19184 12166
rect 19212 12138 19236 12166
rect 19264 12138 19288 12166
rect 19316 12138 19321 12166
rect 2883 11746 2888 11774
rect 2916 11746 2940 11774
rect 2968 11746 2992 11774
rect 3020 11746 3044 11774
rect 3072 11746 3096 11774
rect 3124 11746 3148 11774
rect 3176 11746 3181 11774
rect 20883 11746 20888 11774
rect 20916 11746 20940 11774
rect 20968 11746 20992 11774
rect 21020 11746 21044 11774
rect 21072 11746 21096 11774
rect 21124 11746 21148 11774
rect 21176 11746 21181 11774
rect 1023 11354 1028 11382
rect 1056 11354 1080 11382
rect 1108 11354 1132 11382
rect 1160 11354 1184 11382
rect 1212 11354 1236 11382
rect 1264 11354 1288 11382
rect 1316 11354 1321 11382
rect 19023 11354 19028 11382
rect 19056 11354 19080 11382
rect 19108 11354 19132 11382
rect 19160 11354 19184 11382
rect 19212 11354 19236 11382
rect 19264 11354 19288 11382
rect 19316 11354 19321 11382
rect 2883 10962 2888 10990
rect 2916 10962 2940 10990
rect 2968 10962 2992 10990
rect 3020 10962 3044 10990
rect 3072 10962 3096 10990
rect 3124 10962 3148 10990
rect 3176 10962 3181 10990
rect 20883 10962 20888 10990
rect 20916 10962 20940 10990
rect 20968 10962 20992 10990
rect 21020 10962 21044 10990
rect 21072 10962 21096 10990
rect 21124 10962 21148 10990
rect 21176 10962 21181 10990
rect 1023 10570 1028 10598
rect 1056 10570 1080 10598
rect 1108 10570 1132 10598
rect 1160 10570 1184 10598
rect 1212 10570 1236 10598
rect 1264 10570 1288 10598
rect 1316 10570 1321 10598
rect 19023 10570 19028 10598
rect 19056 10570 19080 10598
rect 19108 10570 19132 10598
rect 19160 10570 19184 10598
rect 19212 10570 19236 10598
rect 19264 10570 19288 10598
rect 19316 10570 19321 10598
rect 2883 10178 2888 10206
rect 2916 10178 2940 10206
rect 2968 10178 2992 10206
rect 3020 10178 3044 10206
rect 3072 10178 3096 10206
rect 3124 10178 3148 10206
rect 3176 10178 3181 10206
rect 20883 10178 20888 10206
rect 20916 10178 20940 10206
rect 20968 10178 20992 10206
rect 21020 10178 21044 10206
rect 21072 10178 21096 10206
rect 21124 10178 21148 10206
rect 21176 10178 21181 10206
rect 1023 9786 1028 9814
rect 1056 9786 1080 9814
rect 1108 9786 1132 9814
rect 1160 9786 1184 9814
rect 1212 9786 1236 9814
rect 1264 9786 1288 9814
rect 1316 9786 1321 9814
rect 19023 9786 19028 9814
rect 19056 9786 19080 9814
rect 19108 9786 19132 9814
rect 19160 9786 19184 9814
rect 19212 9786 19236 9814
rect 19264 9786 19288 9814
rect 19316 9786 19321 9814
rect 2883 9394 2888 9422
rect 2916 9394 2940 9422
rect 2968 9394 2992 9422
rect 3020 9394 3044 9422
rect 3072 9394 3096 9422
rect 3124 9394 3148 9422
rect 3176 9394 3181 9422
rect 20883 9394 20888 9422
rect 20916 9394 20940 9422
rect 20968 9394 20992 9422
rect 21020 9394 21044 9422
rect 21072 9394 21096 9422
rect 21124 9394 21148 9422
rect 21176 9394 21181 9422
rect 1023 9002 1028 9030
rect 1056 9002 1080 9030
rect 1108 9002 1132 9030
rect 1160 9002 1184 9030
rect 1212 9002 1236 9030
rect 1264 9002 1288 9030
rect 1316 9002 1321 9030
rect 19023 9002 19028 9030
rect 19056 9002 19080 9030
rect 19108 9002 19132 9030
rect 19160 9002 19184 9030
rect 19212 9002 19236 9030
rect 19264 9002 19288 9030
rect 19316 9002 19321 9030
rect 2883 8610 2888 8638
rect 2916 8610 2940 8638
rect 2968 8610 2992 8638
rect 3020 8610 3044 8638
rect 3072 8610 3096 8638
rect 3124 8610 3148 8638
rect 3176 8610 3181 8638
rect 20883 8610 20888 8638
rect 20916 8610 20940 8638
rect 20968 8610 20992 8638
rect 21020 8610 21044 8638
rect 21072 8610 21096 8638
rect 21124 8610 21148 8638
rect 21176 8610 21181 8638
rect 1023 8218 1028 8246
rect 1056 8218 1080 8246
rect 1108 8218 1132 8246
rect 1160 8218 1184 8246
rect 1212 8218 1236 8246
rect 1264 8218 1288 8246
rect 1316 8218 1321 8246
rect 19023 8218 19028 8246
rect 19056 8218 19080 8246
rect 19108 8218 19132 8246
rect 19160 8218 19184 8246
rect 19212 8218 19236 8246
rect 19264 8218 19288 8246
rect 19316 8218 19321 8246
rect 2883 7826 2888 7854
rect 2916 7826 2940 7854
rect 2968 7826 2992 7854
rect 3020 7826 3044 7854
rect 3072 7826 3096 7854
rect 3124 7826 3148 7854
rect 3176 7826 3181 7854
rect 20883 7826 20888 7854
rect 20916 7826 20940 7854
rect 20968 7826 20992 7854
rect 21020 7826 21044 7854
rect 21072 7826 21096 7854
rect 21124 7826 21148 7854
rect 21176 7826 21181 7854
rect 1023 7434 1028 7462
rect 1056 7434 1080 7462
rect 1108 7434 1132 7462
rect 1160 7434 1184 7462
rect 1212 7434 1236 7462
rect 1264 7434 1288 7462
rect 1316 7434 1321 7462
rect 19023 7434 19028 7462
rect 19056 7434 19080 7462
rect 19108 7434 19132 7462
rect 19160 7434 19184 7462
rect 19212 7434 19236 7462
rect 19264 7434 19288 7462
rect 19316 7434 19321 7462
rect 2883 7042 2888 7070
rect 2916 7042 2940 7070
rect 2968 7042 2992 7070
rect 3020 7042 3044 7070
rect 3072 7042 3096 7070
rect 3124 7042 3148 7070
rect 3176 7042 3181 7070
rect 20883 7042 20888 7070
rect 20916 7042 20940 7070
rect 20968 7042 20992 7070
rect 21020 7042 21044 7070
rect 21072 7042 21096 7070
rect 21124 7042 21148 7070
rect 21176 7042 21181 7070
rect 1023 6650 1028 6678
rect 1056 6650 1080 6678
rect 1108 6650 1132 6678
rect 1160 6650 1184 6678
rect 1212 6650 1236 6678
rect 1264 6650 1288 6678
rect 1316 6650 1321 6678
rect 19023 6650 19028 6678
rect 19056 6650 19080 6678
rect 19108 6650 19132 6678
rect 19160 6650 19184 6678
rect 19212 6650 19236 6678
rect 19264 6650 19288 6678
rect 19316 6650 19321 6678
rect 2883 6258 2888 6286
rect 2916 6258 2940 6286
rect 2968 6258 2992 6286
rect 3020 6258 3044 6286
rect 3072 6258 3096 6286
rect 3124 6258 3148 6286
rect 3176 6258 3181 6286
rect 20883 6258 20888 6286
rect 20916 6258 20940 6286
rect 20968 6258 20992 6286
rect 21020 6258 21044 6286
rect 21072 6258 21096 6286
rect 21124 6258 21148 6286
rect 21176 6258 21181 6286
rect 14289 6062 14294 6090
rect 14322 6062 16030 6090
rect 16058 6062 16254 6090
rect 16282 6062 16287 6090
rect 12889 6006 12894 6034
rect 12922 6006 13510 6034
rect 13538 6006 13543 6034
rect 1023 5866 1028 5894
rect 1056 5866 1080 5894
rect 1108 5866 1132 5894
rect 1160 5866 1184 5894
rect 1212 5866 1236 5894
rect 1264 5866 1288 5894
rect 1316 5866 1321 5894
rect 19023 5866 19028 5894
rect 19056 5866 19080 5894
rect 19108 5866 19132 5894
rect 19160 5866 19184 5894
rect 19212 5866 19236 5894
rect 19264 5866 19288 5894
rect 19316 5866 19321 5894
rect 12497 5558 12502 5586
rect 12530 5558 13230 5586
rect 13258 5558 22246 5586
rect 22274 5558 22279 5586
rect 2883 5474 2888 5502
rect 2916 5474 2940 5502
rect 2968 5474 2992 5502
rect 3020 5474 3044 5502
rect 3072 5474 3096 5502
rect 3124 5474 3148 5502
rect 3176 5474 3181 5502
rect 20883 5474 20888 5502
rect 20916 5474 20940 5502
rect 20968 5474 20992 5502
rect 21020 5474 21044 5502
rect 21072 5474 21096 5502
rect 21124 5474 21148 5502
rect 21176 5474 21181 5502
rect 6281 5222 6286 5250
rect 6314 5222 12502 5250
rect 12530 5222 12838 5250
rect 12866 5222 12871 5250
rect 12441 5166 12446 5194
rect 12474 5166 14294 5194
rect 14322 5166 14327 5194
rect 1023 5082 1028 5110
rect 1056 5082 1080 5110
rect 1108 5082 1132 5110
rect 1160 5082 1184 5110
rect 1212 5082 1236 5110
rect 1264 5082 1288 5110
rect 1316 5082 1321 5110
rect 19023 5082 19028 5110
rect 19056 5082 19080 5110
rect 19108 5082 19132 5110
rect 19160 5082 19184 5110
rect 19212 5082 19236 5110
rect 19264 5082 19288 5110
rect 19316 5082 19321 5110
rect 10873 4886 10878 4914
rect 10906 4886 11886 4914
rect 11914 4886 11919 4914
rect 12273 4774 12278 4802
rect 12306 4774 13566 4802
rect 13594 4774 18830 4802
rect 18858 4774 18863 4802
rect 2883 4690 2888 4718
rect 2916 4690 2940 4718
rect 2968 4690 2992 4718
rect 3020 4690 3044 4718
rect 3072 4690 3096 4718
rect 3124 4690 3148 4718
rect 3176 4690 3181 4718
rect 20883 4690 20888 4718
rect 20916 4690 20940 4718
rect 20968 4690 20992 4718
rect 21020 4690 21044 4718
rect 21072 4690 21096 4718
rect 21124 4690 21148 4718
rect 21176 4690 21181 4718
rect 1073 4494 1078 4522
rect 1106 4494 1358 4522
rect 1386 4494 11718 4522
rect 11746 4494 11751 4522
rect 1023 4298 1028 4326
rect 1056 4298 1080 4326
rect 1108 4298 1132 4326
rect 1160 4298 1184 4326
rect 1212 4298 1236 4326
rect 1264 4298 1288 4326
rect 1316 4298 1321 4326
rect 19023 4298 19028 4326
rect 19056 4298 19080 4326
rect 19108 4298 19132 4326
rect 19160 4298 19184 4326
rect 19212 4298 19236 4326
rect 19264 4298 19288 4326
rect 19316 4298 19321 4326
rect -480 4186 240 4228
rect -480 4158 910 4186
rect 938 4158 943 4186
rect -480 4116 240 4158
rect 2883 3906 2888 3934
rect 2916 3906 2940 3934
rect 2968 3906 2992 3934
rect 3020 3906 3044 3934
rect 3072 3906 3096 3934
rect 3124 3906 3148 3934
rect 3176 3906 3181 3934
rect 20883 3906 20888 3934
rect 20916 3906 20940 3934
rect 20968 3906 20992 3934
rect 21020 3906 21044 3934
rect 21072 3906 21096 3934
rect 21124 3906 21148 3934
rect 21176 3906 21181 3934
rect 1023 3514 1028 3542
rect 1056 3514 1080 3542
rect 1108 3514 1132 3542
rect 1160 3514 1184 3542
rect 1212 3514 1236 3542
rect 1264 3514 1288 3542
rect 1316 3514 1321 3542
rect 19023 3514 19028 3542
rect 19056 3514 19080 3542
rect 19108 3514 19132 3542
rect 19160 3514 19184 3542
rect 19212 3514 19236 3542
rect 19264 3514 19288 3542
rect 19316 3514 19321 3542
rect 2883 3122 2888 3150
rect 2916 3122 2940 3150
rect 2968 3122 2992 3150
rect 3020 3122 3044 3150
rect 3072 3122 3096 3150
rect 3124 3122 3148 3150
rect 3176 3122 3181 3150
rect 20883 3122 20888 3150
rect 20916 3122 20940 3150
rect 20968 3122 20992 3150
rect 21020 3122 21044 3150
rect 21072 3122 21096 3150
rect 21124 3122 21148 3150
rect 21176 3122 21181 3150
rect 1023 2730 1028 2758
rect 1056 2730 1080 2758
rect 1108 2730 1132 2758
rect 1160 2730 1184 2758
rect 1212 2730 1236 2758
rect 1264 2730 1288 2758
rect 1316 2730 1321 2758
rect 19023 2730 19028 2758
rect 19056 2730 19080 2758
rect 19108 2730 19132 2758
rect 19160 2730 19184 2758
rect 19212 2730 19236 2758
rect 19264 2730 19288 2758
rect 19316 2730 19321 2758
rect 2883 2338 2888 2366
rect 2916 2338 2940 2366
rect 2968 2338 2992 2366
rect 3020 2338 3044 2366
rect 3072 2338 3096 2366
rect 3124 2338 3148 2366
rect 3176 2338 3181 2366
rect 20883 2338 20888 2366
rect 20916 2338 20940 2366
rect 20968 2338 20992 2366
rect 21020 2338 21044 2366
rect 21072 2338 21096 2366
rect 21124 2338 21148 2366
rect 21176 2338 21181 2366
rect 1023 1946 1028 1974
rect 1056 1946 1080 1974
rect 1108 1946 1132 1974
rect 1160 1946 1184 1974
rect 1212 1946 1236 1974
rect 1264 1946 1288 1974
rect 1316 1946 1321 1974
rect 19023 1946 19028 1974
rect 19056 1946 19080 1974
rect 19108 1946 19132 1974
rect 19160 1946 19184 1974
rect 19212 1946 19236 1974
rect 19264 1946 19288 1974
rect 19316 1946 19321 1974
rect 18657 1694 18662 1722
rect 18690 1694 18998 1722
rect 19026 1694 19031 1722
rect 2883 1554 2888 1582
rect 2916 1554 2940 1582
rect 2968 1554 2992 1582
rect 3020 1554 3044 1582
rect 3072 1554 3096 1582
rect 3124 1554 3148 1582
rect 3176 1554 3181 1582
rect 20883 1554 20888 1582
rect 20916 1554 20940 1582
rect 20968 1554 20992 1582
rect 21020 1554 21044 1582
rect 21072 1554 21096 1582
rect 21124 1554 21148 1582
rect 21176 1554 21181 1582
<< via3 >>
rect 1028 23114 1056 23142
rect 1080 23114 1108 23142
rect 1132 23114 1160 23142
rect 1184 23114 1212 23142
rect 1236 23114 1264 23142
rect 1288 23114 1316 23142
rect 19028 23114 19056 23142
rect 19080 23114 19108 23142
rect 19132 23114 19160 23142
rect 19184 23114 19212 23142
rect 19236 23114 19264 23142
rect 19288 23114 19316 23142
rect 2888 22722 2916 22750
rect 2940 22722 2968 22750
rect 2992 22722 3020 22750
rect 3044 22722 3072 22750
rect 3096 22722 3124 22750
rect 3148 22722 3176 22750
rect 20888 22722 20916 22750
rect 20940 22722 20968 22750
rect 20992 22722 21020 22750
rect 21044 22722 21072 22750
rect 21096 22722 21124 22750
rect 21148 22722 21176 22750
rect 1028 22330 1056 22358
rect 1080 22330 1108 22358
rect 1132 22330 1160 22358
rect 1184 22330 1212 22358
rect 1236 22330 1264 22358
rect 1288 22330 1316 22358
rect 19028 22330 19056 22358
rect 19080 22330 19108 22358
rect 19132 22330 19160 22358
rect 19184 22330 19212 22358
rect 19236 22330 19264 22358
rect 19288 22330 19316 22358
rect 2888 21938 2916 21966
rect 2940 21938 2968 21966
rect 2992 21938 3020 21966
rect 3044 21938 3072 21966
rect 3096 21938 3124 21966
rect 3148 21938 3176 21966
rect 20888 21938 20916 21966
rect 20940 21938 20968 21966
rect 20992 21938 21020 21966
rect 21044 21938 21072 21966
rect 21096 21938 21124 21966
rect 21148 21938 21176 21966
rect 1028 21546 1056 21574
rect 1080 21546 1108 21574
rect 1132 21546 1160 21574
rect 1184 21546 1212 21574
rect 1236 21546 1264 21574
rect 1288 21546 1316 21574
rect 19028 21546 19056 21574
rect 19080 21546 19108 21574
rect 19132 21546 19160 21574
rect 19184 21546 19212 21574
rect 19236 21546 19264 21574
rect 19288 21546 19316 21574
rect 2888 21154 2916 21182
rect 2940 21154 2968 21182
rect 2992 21154 3020 21182
rect 3044 21154 3072 21182
rect 3096 21154 3124 21182
rect 3148 21154 3176 21182
rect 20888 21154 20916 21182
rect 20940 21154 20968 21182
rect 20992 21154 21020 21182
rect 21044 21154 21072 21182
rect 21096 21154 21124 21182
rect 21148 21154 21176 21182
rect 1028 20762 1056 20790
rect 1080 20762 1108 20790
rect 1132 20762 1160 20790
rect 1184 20762 1212 20790
rect 1236 20762 1264 20790
rect 1288 20762 1316 20790
rect 19028 20762 19056 20790
rect 19080 20762 19108 20790
rect 19132 20762 19160 20790
rect 19184 20762 19212 20790
rect 19236 20762 19264 20790
rect 19288 20762 19316 20790
rect 2888 20370 2916 20398
rect 2940 20370 2968 20398
rect 2992 20370 3020 20398
rect 3044 20370 3072 20398
rect 3096 20370 3124 20398
rect 3148 20370 3176 20398
rect 20888 20370 20916 20398
rect 20940 20370 20968 20398
rect 20992 20370 21020 20398
rect 21044 20370 21072 20398
rect 21096 20370 21124 20398
rect 21148 20370 21176 20398
rect 1028 19978 1056 20006
rect 1080 19978 1108 20006
rect 1132 19978 1160 20006
rect 1184 19978 1212 20006
rect 1236 19978 1264 20006
rect 1288 19978 1316 20006
rect 19028 19978 19056 20006
rect 19080 19978 19108 20006
rect 19132 19978 19160 20006
rect 19184 19978 19212 20006
rect 19236 19978 19264 20006
rect 19288 19978 19316 20006
rect 2888 19586 2916 19614
rect 2940 19586 2968 19614
rect 2992 19586 3020 19614
rect 3044 19586 3072 19614
rect 3096 19586 3124 19614
rect 3148 19586 3176 19614
rect 20888 19586 20916 19614
rect 20940 19586 20968 19614
rect 20992 19586 21020 19614
rect 21044 19586 21072 19614
rect 21096 19586 21124 19614
rect 21148 19586 21176 19614
rect 1028 19194 1056 19222
rect 1080 19194 1108 19222
rect 1132 19194 1160 19222
rect 1184 19194 1212 19222
rect 1236 19194 1264 19222
rect 1288 19194 1316 19222
rect 19028 19194 19056 19222
rect 19080 19194 19108 19222
rect 19132 19194 19160 19222
rect 19184 19194 19212 19222
rect 19236 19194 19264 19222
rect 19288 19194 19316 19222
rect 2888 18802 2916 18830
rect 2940 18802 2968 18830
rect 2992 18802 3020 18830
rect 3044 18802 3072 18830
rect 3096 18802 3124 18830
rect 3148 18802 3176 18830
rect 20888 18802 20916 18830
rect 20940 18802 20968 18830
rect 20992 18802 21020 18830
rect 21044 18802 21072 18830
rect 21096 18802 21124 18830
rect 21148 18802 21176 18830
rect 1028 18410 1056 18438
rect 1080 18410 1108 18438
rect 1132 18410 1160 18438
rect 1184 18410 1212 18438
rect 1236 18410 1264 18438
rect 1288 18410 1316 18438
rect 19028 18410 19056 18438
rect 19080 18410 19108 18438
rect 19132 18410 19160 18438
rect 19184 18410 19212 18438
rect 19236 18410 19264 18438
rect 19288 18410 19316 18438
rect 2888 18018 2916 18046
rect 2940 18018 2968 18046
rect 2992 18018 3020 18046
rect 3044 18018 3072 18046
rect 3096 18018 3124 18046
rect 3148 18018 3176 18046
rect 20888 18018 20916 18046
rect 20940 18018 20968 18046
rect 20992 18018 21020 18046
rect 21044 18018 21072 18046
rect 21096 18018 21124 18046
rect 21148 18018 21176 18046
rect 1028 17626 1056 17654
rect 1080 17626 1108 17654
rect 1132 17626 1160 17654
rect 1184 17626 1212 17654
rect 1236 17626 1264 17654
rect 1288 17626 1316 17654
rect 19028 17626 19056 17654
rect 19080 17626 19108 17654
rect 19132 17626 19160 17654
rect 19184 17626 19212 17654
rect 19236 17626 19264 17654
rect 19288 17626 19316 17654
rect 2888 17234 2916 17262
rect 2940 17234 2968 17262
rect 2992 17234 3020 17262
rect 3044 17234 3072 17262
rect 3096 17234 3124 17262
rect 3148 17234 3176 17262
rect 20888 17234 20916 17262
rect 20940 17234 20968 17262
rect 20992 17234 21020 17262
rect 21044 17234 21072 17262
rect 21096 17234 21124 17262
rect 21148 17234 21176 17262
rect 1028 16842 1056 16870
rect 1080 16842 1108 16870
rect 1132 16842 1160 16870
rect 1184 16842 1212 16870
rect 1236 16842 1264 16870
rect 1288 16842 1316 16870
rect 19028 16842 19056 16870
rect 19080 16842 19108 16870
rect 19132 16842 19160 16870
rect 19184 16842 19212 16870
rect 19236 16842 19264 16870
rect 19288 16842 19316 16870
rect 2888 16450 2916 16478
rect 2940 16450 2968 16478
rect 2992 16450 3020 16478
rect 3044 16450 3072 16478
rect 3096 16450 3124 16478
rect 3148 16450 3176 16478
rect 20888 16450 20916 16478
rect 20940 16450 20968 16478
rect 20992 16450 21020 16478
rect 21044 16450 21072 16478
rect 21096 16450 21124 16478
rect 21148 16450 21176 16478
rect 1028 16058 1056 16086
rect 1080 16058 1108 16086
rect 1132 16058 1160 16086
rect 1184 16058 1212 16086
rect 1236 16058 1264 16086
rect 1288 16058 1316 16086
rect 19028 16058 19056 16086
rect 19080 16058 19108 16086
rect 19132 16058 19160 16086
rect 19184 16058 19212 16086
rect 19236 16058 19264 16086
rect 19288 16058 19316 16086
rect 2888 15666 2916 15694
rect 2940 15666 2968 15694
rect 2992 15666 3020 15694
rect 3044 15666 3072 15694
rect 3096 15666 3124 15694
rect 3148 15666 3176 15694
rect 20888 15666 20916 15694
rect 20940 15666 20968 15694
rect 20992 15666 21020 15694
rect 21044 15666 21072 15694
rect 21096 15666 21124 15694
rect 21148 15666 21176 15694
rect 1028 15274 1056 15302
rect 1080 15274 1108 15302
rect 1132 15274 1160 15302
rect 1184 15274 1212 15302
rect 1236 15274 1264 15302
rect 1288 15274 1316 15302
rect 19028 15274 19056 15302
rect 19080 15274 19108 15302
rect 19132 15274 19160 15302
rect 19184 15274 19212 15302
rect 19236 15274 19264 15302
rect 19288 15274 19316 15302
rect 2888 14882 2916 14910
rect 2940 14882 2968 14910
rect 2992 14882 3020 14910
rect 3044 14882 3072 14910
rect 3096 14882 3124 14910
rect 3148 14882 3176 14910
rect 20888 14882 20916 14910
rect 20940 14882 20968 14910
rect 20992 14882 21020 14910
rect 21044 14882 21072 14910
rect 21096 14882 21124 14910
rect 21148 14882 21176 14910
rect 1028 14490 1056 14518
rect 1080 14490 1108 14518
rect 1132 14490 1160 14518
rect 1184 14490 1212 14518
rect 1236 14490 1264 14518
rect 1288 14490 1316 14518
rect 19028 14490 19056 14518
rect 19080 14490 19108 14518
rect 19132 14490 19160 14518
rect 19184 14490 19212 14518
rect 19236 14490 19264 14518
rect 19288 14490 19316 14518
rect 2888 14098 2916 14126
rect 2940 14098 2968 14126
rect 2992 14098 3020 14126
rect 3044 14098 3072 14126
rect 3096 14098 3124 14126
rect 3148 14098 3176 14126
rect 20888 14098 20916 14126
rect 20940 14098 20968 14126
rect 20992 14098 21020 14126
rect 21044 14098 21072 14126
rect 21096 14098 21124 14126
rect 21148 14098 21176 14126
rect 1028 13706 1056 13734
rect 1080 13706 1108 13734
rect 1132 13706 1160 13734
rect 1184 13706 1212 13734
rect 1236 13706 1264 13734
rect 1288 13706 1316 13734
rect 19028 13706 19056 13734
rect 19080 13706 19108 13734
rect 19132 13706 19160 13734
rect 19184 13706 19212 13734
rect 19236 13706 19264 13734
rect 19288 13706 19316 13734
rect 2888 13314 2916 13342
rect 2940 13314 2968 13342
rect 2992 13314 3020 13342
rect 3044 13314 3072 13342
rect 3096 13314 3124 13342
rect 3148 13314 3176 13342
rect 20888 13314 20916 13342
rect 20940 13314 20968 13342
rect 20992 13314 21020 13342
rect 21044 13314 21072 13342
rect 21096 13314 21124 13342
rect 21148 13314 21176 13342
rect 1028 12922 1056 12950
rect 1080 12922 1108 12950
rect 1132 12922 1160 12950
rect 1184 12922 1212 12950
rect 1236 12922 1264 12950
rect 1288 12922 1316 12950
rect 19028 12922 19056 12950
rect 19080 12922 19108 12950
rect 19132 12922 19160 12950
rect 19184 12922 19212 12950
rect 19236 12922 19264 12950
rect 19288 12922 19316 12950
rect 2888 12530 2916 12558
rect 2940 12530 2968 12558
rect 2992 12530 3020 12558
rect 3044 12530 3072 12558
rect 3096 12530 3124 12558
rect 3148 12530 3176 12558
rect 20888 12530 20916 12558
rect 20940 12530 20968 12558
rect 20992 12530 21020 12558
rect 21044 12530 21072 12558
rect 21096 12530 21124 12558
rect 21148 12530 21176 12558
rect 1028 12138 1056 12166
rect 1080 12138 1108 12166
rect 1132 12138 1160 12166
rect 1184 12138 1212 12166
rect 1236 12138 1264 12166
rect 1288 12138 1316 12166
rect 19028 12138 19056 12166
rect 19080 12138 19108 12166
rect 19132 12138 19160 12166
rect 19184 12138 19212 12166
rect 19236 12138 19264 12166
rect 19288 12138 19316 12166
rect 2888 11746 2916 11774
rect 2940 11746 2968 11774
rect 2992 11746 3020 11774
rect 3044 11746 3072 11774
rect 3096 11746 3124 11774
rect 3148 11746 3176 11774
rect 20888 11746 20916 11774
rect 20940 11746 20968 11774
rect 20992 11746 21020 11774
rect 21044 11746 21072 11774
rect 21096 11746 21124 11774
rect 21148 11746 21176 11774
rect 1028 11354 1056 11382
rect 1080 11354 1108 11382
rect 1132 11354 1160 11382
rect 1184 11354 1212 11382
rect 1236 11354 1264 11382
rect 1288 11354 1316 11382
rect 19028 11354 19056 11382
rect 19080 11354 19108 11382
rect 19132 11354 19160 11382
rect 19184 11354 19212 11382
rect 19236 11354 19264 11382
rect 19288 11354 19316 11382
rect 2888 10962 2916 10990
rect 2940 10962 2968 10990
rect 2992 10962 3020 10990
rect 3044 10962 3072 10990
rect 3096 10962 3124 10990
rect 3148 10962 3176 10990
rect 20888 10962 20916 10990
rect 20940 10962 20968 10990
rect 20992 10962 21020 10990
rect 21044 10962 21072 10990
rect 21096 10962 21124 10990
rect 21148 10962 21176 10990
rect 1028 10570 1056 10598
rect 1080 10570 1108 10598
rect 1132 10570 1160 10598
rect 1184 10570 1212 10598
rect 1236 10570 1264 10598
rect 1288 10570 1316 10598
rect 19028 10570 19056 10598
rect 19080 10570 19108 10598
rect 19132 10570 19160 10598
rect 19184 10570 19212 10598
rect 19236 10570 19264 10598
rect 19288 10570 19316 10598
rect 2888 10178 2916 10206
rect 2940 10178 2968 10206
rect 2992 10178 3020 10206
rect 3044 10178 3072 10206
rect 3096 10178 3124 10206
rect 3148 10178 3176 10206
rect 20888 10178 20916 10206
rect 20940 10178 20968 10206
rect 20992 10178 21020 10206
rect 21044 10178 21072 10206
rect 21096 10178 21124 10206
rect 21148 10178 21176 10206
rect 1028 9786 1056 9814
rect 1080 9786 1108 9814
rect 1132 9786 1160 9814
rect 1184 9786 1212 9814
rect 1236 9786 1264 9814
rect 1288 9786 1316 9814
rect 19028 9786 19056 9814
rect 19080 9786 19108 9814
rect 19132 9786 19160 9814
rect 19184 9786 19212 9814
rect 19236 9786 19264 9814
rect 19288 9786 19316 9814
rect 2888 9394 2916 9422
rect 2940 9394 2968 9422
rect 2992 9394 3020 9422
rect 3044 9394 3072 9422
rect 3096 9394 3124 9422
rect 3148 9394 3176 9422
rect 20888 9394 20916 9422
rect 20940 9394 20968 9422
rect 20992 9394 21020 9422
rect 21044 9394 21072 9422
rect 21096 9394 21124 9422
rect 21148 9394 21176 9422
rect 1028 9002 1056 9030
rect 1080 9002 1108 9030
rect 1132 9002 1160 9030
rect 1184 9002 1212 9030
rect 1236 9002 1264 9030
rect 1288 9002 1316 9030
rect 19028 9002 19056 9030
rect 19080 9002 19108 9030
rect 19132 9002 19160 9030
rect 19184 9002 19212 9030
rect 19236 9002 19264 9030
rect 19288 9002 19316 9030
rect 2888 8610 2916 8638
rect 2940 8610 2968 8638
rect 2992 8610 3020 8638
rect 3044 8610 3072 8638
rect 3096 8610 3124 8638
rect 3148 8610 3176 8638
rect 20888 8610 20916 8638
rect 20940 8610 20968 8638
rect 20992 8610 21020 8638
rect 21044 8610 21072 8638
rect 21096 8610 21124 8638
rect 21148 8610 21176 8638
rect 1028 8218 1056 8246
rect 1080 8218 1108 8246
rect 1132 8218 1160 8246
rect 1184 8218 1212 8246
rect 1236 8218 1264 8246
rect 1288 8218 1316 8246
rect 19028 8218 19056 8246
rect 19080 8218 19108 8246
rect 19132 8218 19160 8246
rect 19184 8218 19212 8246
rect 19236 8218 19264 8246
rect 19288 8218 19316 8246
rect 2888 7826 2916 7854
rect 2940 7826 2968 7854
rect 2992 7826 3020 7854
rect 3044 7826 3072 7854
rect 3096 7826 3124 7854
rect 3148 7826 3176 7854
rect 20888 7826 20916 7854
rect 20940 7826 20968 7854
rect 20992 7826 21020 7854
rect 21044 7826 21072 7854
rect 21096 7826 21124 7854
rect 21148 7826 21176 7854
rect 1028 7434 1056 7462
rect 1080 7434 1108 7462
rect 1132 7434 1160 7462
rect 1184 7434 1212 7462
rect 1236 7434 1264 7462
rect 1288 7434 1316 7462
rect 19028 7434 19056 7462
rect 19080 7434 19108 7462
rect 19132 7434 19160 7462
rect 19184 7434 19212 7462
rect 19236 7434 19264 7462
rect 19288 7434 19316 7462
rect 2888 7042 2916 7070
rect 2940 7042 2968 7070
rect 2992 7042 3020 7070
rect 3044 7042 3072 7070
rect 3096 7042 3124 7070
rect 3148 7042 3176 7070
rect 20888 7042 20916 7070
rect 20940 7042 20968 7070
rect 20992 7042 21020 7070
rect 21044 7042 21072 7070
rect 21096 7042 21124 7070
rect 21148 7042 21176 7070
rect 1028 6650 1056 6678
rect 1080 6650 1108 6678
rect 1132 6650 1160 6678
rect 1184 6650 1212 6678
rect 1236 6650 1264 6678
rect 1288 6650 1316 6678
rect 19028 6650 19056 6678
rect 19080 6650 19108 6678
rect 19132 6650 19160 6678
rect 19184 6650 19212 6678
rect 19236 6650 19264 6678
rect 19288 6650 19316 6678
rect 2888 6258 2916 6286
rect 2940 6258 2968 6286
rect 2992 6258 3020 6286
rect 3044 6258 3072 6286
rect 3096 6258 3124 6286
rect 3148 6258 3176 6286
rect 20888 6258 20916 6286
rect 20940 6258 20968 6286
rect 20992 6258 21020 6286
rect 21044 6258 21072 6286
rect 21096 6258 21124 6286
rect 21148 6258 21176 6286
rect 1028 5866 1056 5894
rect 1080 5866 1108 5894
rect 1132 5866 1160 5894
rect 1184 5866 1212 5894
rect 1236 5866 1264 5894
rect 1288 5866 1316 5894
rect 19028 5866 19056 5894
rect 19080 5866 19108 5894
rect 19132 5866 19160 5894
rect 19184 5866 19212 5894
rect 19236 5866 19264 5894
rect 19288 5866 19316 5894
rect 2888 5474 2916 5502
rect 2940 5474 2968 5502
rect 2992 5474 3020 5502
rect 3044 5474 3072 5502
rect 3096 5474 3124 5502
rect 3148 5474 3176 5502
rect 20888 5474 20916 5502
rect 20940 5474 20968 5502
rect 20992 5474 21020 5502
rect 21044 5474 21072 5502
rect 21096 5474 21124 5502
rect 21148 5474 21176 5502
rect 1028 5082 1056 5110
rect 1080 5082 1108 5110
rect 1132 5082 1160 5110
rect 1184 5082 1212 5110
rect 1236 5082 1264 5110
rect 1288 5082 1316 5110
rect 19028 5082 19056 5110
rect 19080 5082 19108 5110
rect 19132 5082 19160 5110
rect 19184 5082 19212 5110
rect 19236 5082 19264 5110
rect 19288 5082 19316 5110
rect 2888 4690 2916 4718
rect 2940 4690 2968 4718
rect 2992 4690 3020 4718
rect 3044 4690 3072 4718
rect 3096 4690 3124 4718
rect 3148 4690 3176 4718
rect 20888 4690 20916 4718
rect 20940 4690 20968 4718
rect 20992 4690 21020 4718
rect 21044 4690 21072 4718
rect 21096 4690 21124 4718
rect 21148 4690 21176 4718
rect 1028 4298 1056 4326
rect 1080 4298 1108 4326
rect 1132 4298 1160 4326
rect 1184 4298 1212 4326
rect 1236 4298 1264 4326
rect 1288 4298 1316 4326
rect 19028 4298 19056 4326
rect 19080 4298 19108 4326
rect 19132 4298 19160 4326
rect 19184 4298 19212 4326
rect 19236 4298 19264 4326
rect 19288 4298 19316 4326
rect 2888 3906 2916 3934
rect 2940 3906 2968 3934
rect 2992 3906 3020 3934
rect 3044 3906 3072 3934
rect 3096 3906 3124 3934
rect 3148 3906 3176 3934
rect 20888 3906 20916 3934
rect 20940 3906 20968 3934
rect 20992 3906 21020 3934
rect 21044 3906 21072 3934
rect 21096 3906 21124 3934
rect 21148 3906 21176 3934
rect 1028 3514 1056 3542
rect 1080 3514 1108 3542
rect 1132 3514 1160 3542
rect 1184 3514 1212 3542
rect 1236 3514 1264 3542
rect 1288 3514 1316 3542
rect 19028 3514 19056 3542
rect 19080 3514 19108 3542
rect 19132 3514 19160 3542
rect 19184 3514 19212 3542
rect 19236 3514 19264 3542
rect 19288 3514 19316 3542
rect 2888 3122 2916 3150
rect 2940 3122 2968 3150
rect 2992 3122 3020 3150
rect 3044 3122 3072 3150
rect 3096 3122 3124 3150
rect 3148 3122 3176 3150
rect 20888 3122 20916 3150
rect 20940 3122 20968 3150
rect 20992 3122 21020 3150
rect 21044 3122 21072 3150
rect 21096 3122 21124 3150
rect 21148 3122 21176 3150
rect 1028 2730 1056 2758
rect 1080 2730 1108 2758
rect 1132 2730 1160 2758
rect 1184 2730 1212 2758
rect 1236 2730 1264 2758
rect 1288 2730 1316 2758
rect 19028 2730 19056 2758
rect 19080 2730 19108 2758
rect 19132 2730 19160 2758
rect 19184 2730 19212 2758
rect 19236 2730 19264 2758
rect 19288 2730 19316 2758
rect 2888 2338 2916 2366
rect 2940 2338 2968 2366
rect 2992 2338 3020 2366
rect 3044 2338 3072 2366
rect 3096 2338 3124 2366
rect 3148 2338 3176 2366
rect 20888 2338 20916 2366
rect 20940 2338 20968 2366
rect 20992 2338 21020 2366
rect 21044 2338 21072 2366
rect 21096 2338 21124 2366
rect 21148 2338 21176 2366
rect 1028 1946 1056 1974
rect 1080 1946 1108 1974
rect 1132 1946 1160 1974
rect 1184 1946 1212 1974
rect 1236 1946 1264 1974
rect 1288 1946 1316 1974
rect 19028 1946 19056 1974
rect 19080 1946 19108 1974
rect 19132 1946 19160 1974
rect 19184 1946 19212 1974
rect 19236 1946 19264 1974
rect 19288 1946 19316 1974
rect 2888 1554 2916 1582
rect 2940 1554 2968 1582
rect 2992 1554 3020 1582
rect 3044 1554 3072 1582
rect 3096 1554 3124 1582
rect 3148 1554 3176 1582
rect 20888 1554 20916 1582
rect 20940 1554 20968 1582
rect 20992 1554 21020 1582
rect 21044 1554 21072 1582
rect 21096 1554 21124 1582
rect 21148 1554 21176 1582
<< metal4 >>
rect 1017 23142 1327 23158
rect 1017 23114 1028 23142
rect 1056 23114 1080 23142
rect 1108 23114 1132 23142
rect 1160 23114 1184 23142
rect 1212 23114 1236 23142
rect 1264 23114 1288 23142
rect 1316 23114 1327 23142
rect 1017 22358 1327 23114
rect 1017 22330 1028 22358
rect 1056 22330 1080 22358
rect 1108 22330 1132 22358
rect 1160 22330 1184 22358
rect 1212 22330 1236 22358
rect 1264 22330 1288 22358
rect 1316 22330 1327 22358
rect 1017 21574 1327 22330
rect 1017 21546 1028 21574
rect 1056 21546 1080 21574
rect 1108 21546 1132 21574
rect 1160 21546 1184 21574
rect 1212 21546 1236 21574
rect 1264 21546 1288 21574
rect 1316 21546 1327 21574
rect 1017 20790 1327 21546
rect 1017 20762 1028 20790
rect 1056 20762 1080 20790
rect 1108 20762 1132 20790
rect 1160 20762 1184 20790
rect 1212 20762 1236 20790
rect 1264 20762 1288 20790
rect 1316 20762 1327 20790
rect 1017 20006 1327 20762
rect 1017 19978 1028 20006
rect 1056 19978 1080 20006
rect 1108 19978 1132 20006
rect 1160 19978 1184 20006
rect 1212 19978 1236 20006
rect 1264 19978 1288 20006
rect 1316 19978 1327 20006
rect 1017 19222 1327 19978
rect 1017 19194 1028 19222
rect 1056 19194 1080 19222
rect 1108 19194 1132 19222
rect 1160 19194 1184 19222
rect 1212 19194 1236 19222
rect 1264 19194 1288 19222
rect 1316 19194 1327 19222
rect 1017 18438 1327 19194
rect 1017 18410 1028 18438
rect 1056 18410 1080 18438
rect 1108 18410 1132 18438
rect 1160 18410 1184 18438
rect 1212 18410 1236 18438
rect 1264 18410 1288 18438
rect 1316 18410 1327 18438
rect 1017 17654 1327 18410
rect 1017 17626 1028 17654
rect 1056 17626 1080 17654
rect 1108 17626 1132 17654
rect 1160 17626 1184 17654
rect 1212 17626 1236 17654
rect 1264 17626 1288 17654
rect 1316 17626 1327 17654
rect 1017 16870 1327 17626
rect 1017 16842 1028 16870
rect 1056 16842 1080 16870
rect 1108 16842 1132 16870
rect 1160 16842 1184 16870
rect 1212 16842 1236 16870
rect 1264 16842 1288 16870
rect 1316 16842 1327 16870
rect 1017 16086 1327 16842
rect 1017 16058 1028 16086
rect 1056 16058 1080 16086
rect 1108 16058 1132 16086
rect 1160 16058 1184 16086
rect 1212 16058 1236 16086
rect 1264 16058 1288 16086
rect 1316 16058 1327 16086
rect 1017 15302 1327 16058
rect 1017 15274 1028 15302
rect 1056 15274 1080 15302
rect 1108 15274 1132 15302
rect 1160 15274 1184 15302
rect 1212 15274 1236 15302
rect 1264 15274 1288 15302
rect 1316 15274 1327 15302
rect 1017 14518 1327 15274
rect 1017 14490 1028 14518
rect 1056 14490 1080 14518
rect 1108 14490 1132 14518
rect 1160 14490 1184 14518
rect 1212 14490 1236 14518
rect 1264 14490 1288 14518
rect 1316 14490 1327 14518
rect 1017 13734 1327 14490
rect 1017 13706 1028 13734
rect 1056 13706 1080 13734
rect 1108 13706 1132 13734
rect 1160 13706 1184 13734
rect 1212 13706 1236 13734
rect 1264 13706 1288 13734
rect 1316 13706 1327 13734
rect 1017 12950 1327 13706
rect 1017 12922 1028 12950
rect 1056 12922 1080 12950
rect 1108 12922 1132 12950
rect 1160 12922 1184 12950
rect 1212 12922 1236 12950
rect 1264 12922 1288 12950
rect 1316 12922 1327 12950
rect 1017 12166 1327 12922
rect 1017 12138 1028 12166
rect 1056 12138 1080 12166
rect 1108 12138 1132 12166
rect 1160 12138 1184 12166
rect 1212 12138 1236 12166
rect 1264 12138 1288 12166
rect 1316 12138 1327 12166
rect 1017 11382 1327 12138
rect 1017 11354 1028 11382
rect 1056 11354 1080 11382
rect 1108 11354 1132 11382
rect 1160 11354 1184 11382
rect 1212 11354 1236 11382
rect 1264 11354 1288 11382
rect 1316 11354 1327 11382
rect 1017 10598 1327 11354
rect 1017 10570 1028 10598
rect 1056 10570 1080 10598
rect 1108 10570 1132 10598
rect 1160 10570 1184 10598
rect 1212 10570 1236 10598
rect 1264 10570 1288 10598
rect 1316 10570 1327 10598
rect 1017 9814 1327 10570
rect 1017 9786 1028 9814
rect 1056 9786 1080 9814
rect 1108 9786 1132 9814
rect 1160 9786 1184 9814
rect 1212 9786 1236 9814
rect 1264 9786 1288 9814
rect 1316 9786 1327 9814
rect 1017 9030 1327 9786
rect 1017 9002 1028 9030
rect 1056 9002 1080 9030
rect 1108 9002 1132 9030
rect 1160 9002 1184 9030
rect 1212 9002 1236 9030
rect 1264 9002 1288 9030
rect 1316 9002 1327 9030
rect 1017 8246 1327 9002
rect 1017 8218 1028 8246
rect 1056 8218 1080 8246
rect 1108 8218 1132 8246
rect 1160 8218 1184 8246
rect 1212 8218 1236 8246
rect 1264 8218 1288 8246
rect 1316 8218 1327 8246
rect 1017 7462 1327 8218
rect 1017 7434 1028 7462
rect 1056 7434 1080 7462
rect 1108 7434 1132 7462
rect 1160 7434 1184 7462
rect 1212 7434 1236 7462
rect 1264 7434 1288 7462
rect 1316 7434 1327 7462
rect 1017 6678 1327 7434
rect 1017 6650 1028 6678
rect 1056 6650 1080 6678
rect 1108 6650 1132 6678
rect 1160 6650 1184 6678
rect 1212 6650 1236 6678
rect 1264 6650 1288 6678
rect 1316 6650 1327 6678
rect 1017 5894 1327 6650
rect 1017 5866 1028 5894
rect 1056 5866 1080 5894
rect 1108 5866 1132 5894
rect 1160 5866 1184 5894
rect 1212 5866 1236 5894
rect 1264 5866 1288 5894
rect 1316 5866 1327 5894
rect 1017 5110 1327 5866
rect 1017 5082 1028 5110
rect 1056 5082 1080 5110
rect 1108 5082 1132 5110
rect 1160 5082 1184 5110
rect 1212 5082 1236 5110
rect 1264 5082 1288 5110
rect 1316 5082 1327 5110
rect 1017 4326 1327 5082
rect 1017 4298 1028 4326
rect 1056 4298 1080 4326
rect 1108 4298 1132 4326
rect 1160 4298 1184 4326
rect 1212 4298 1236 4326
rect 1264 4298 1288 4326
rect 1316 4298 1327 4326
rect 1017 3542 1327 4298
rect 1017 3514 1028 3542
rect 1056 3514 1080 3542
rect 1108 3514 1132 3542
rect 1160 3514 1184 3542
rect 1212 3514 1236 3542
rect 1264 3514 1288 3542
rect 1316 3514 1327 3542
rect 1017 2758 1327 3514
rect 1017 2730 1028 2758
rect 1056 2730 1080 2758
rect 1108 2730 1132 2758
rect 1160 2730 1184 2758
rect 1212 2730 1236 2758
rect 1264 2730 1288 2758
rect 1316 2730 1327 2758
rect 1017 1974 1327 2730
rect 1017 1946 1028 1974
rect 1056 1946 1080 1974
rect 1108 1946 1132 1974
rect 1160 1946 1184 1974
rect 1212 1946 1236 1974
rect 1264 1946 1288 1974
rect 1316 1946 1327 1974
rect 1017 1538 1327 1946
rect 2877 22750 3187 23158
rect 2877 22722 2888 22750
rect 2916 22722 2940 22750
rect 2968 22722 2992 22750
rect 3020 22722 3044 22750
rect 3072 22722 3096 22750
rect 3124 22722 3148 22750
rect 3176 22722 3187 22750
rect 2877 21966 3187 22722
rect 2877 21938 2888 21966
rect 2916 21938 2940 21966
rect 2968 21938 2992 21966
rect 3020 21938 3044 21966
rect 3072 21938 3096 21966
rect 3124 21938 3148 21966
rect 3176 21938 3187 21966
rect 2877 21182 3187 21938
rect 2877 21154 2888 21182
rect 2916 21154 2940 21182
rect 2968 21154 2992 21182
rect 3020 21154 3044 21182
rect 3072 21154 3096 21182
rect 3124 21154 3148 21182
rect 3176 21154 3187 21182
rect 2877 20398 3187 21154
rect 2877 20370 2888 20398
rect 2916 20370 2940 20398
rect 2968 20370 2992 20398
rect 3020 20370 3044 20398
rect 3072 20370 3096 20398
rect 3124 20370 3148 20398
rect 3176 20370 3187 20398
rect 2877 19614 3187 20370
rect 2877 19586 2888 19614
rect 2916 19586 2940 19614
rect 2968 19586 2992 19614
rect 3020 19586 3044 19614
rect 3072 19586 3096 19614
rect 3124 19586 3148 19614
rect 3176 19586 3187 19614
rect 2877 18830 3187 19586
rect 2877 18802 2888 18830
rect 2916 18802 2940 18830
rect 2968 18802 2992 18830
rect 3020 18802 3044 18830
rect 3072 18802 3096 18830
rect 3124 18802 3148 18830
rect 3176 18802 3187 18830
rect 2877 18046 3187 18802
rect 2877 18018 2888 18046
rect 2916 18018 2940 18046
rect 2968 18018 2992 18046
rect 3020 18018 3044 18046
rect 3072 18018 3096 18046
rect 3124 18018 3148 18046
rect 3176 18018 3187 18046
rect 2877 17262 3187 18018
rect 2877 17234 2888 17262
rect 2916 17234 2940 17262
rect 2968 17234 2992 17262
rect 3020 17234 3044 17262
rect 3072 17234 3096 17262
rect 3124 17234 3148 17262
rect 3176 17234 3187 17262
rect 2877 16478 3187 17234
rect 2877 16450 2888 16478
rect 2916 16450 2940 16478
rect 2968 16450 2992 16478
rect 3020 16450 3044 16478
rect 3072 16450 3096 16478
rect 3124 16450 3148 16478
rect 3176 16450 3187 16478
rect 2877 15694 3187 16450
rect 2877 15666 2888 15694
rect 2916 15666 2940 15694
rect 2968 15666 2992 15694
rect 3020 15666 3044 15694
rect 3072 15666 3096 15694
rect 3124 15666 3148 15694
rect 3176 15666 3187 15694
rect 2877 14910 3187 15666
rect 2877 14882 2888 14910
rect 2916 14882 2940 14910
rect 2968 14882 2992 14910
rect 3020 14882 3044 14910
rect 3072 14882 3096 14910
rect 3124 14882 3148 14910
rect 3176 14882 3187 14910
rect 2877 14126 3187 14882
rect 2877 14098 2888 14126
rect 2916 14098 2940 14126
rect 2968 14098 2992 14126
rect 3020 14098 3044 14126
rect 3072 14098 3096 14126
rect 3124 14098 3148 14126
rect 3176 14098 3187 14126
rect 2877 13342 3187 14098
rect 2877 13314 2888 13342
rect 2916 13314 2940 13342
rect 2968 13314 2992 13342
rect 3020 13314 3044 13342
rect 3072 13314 3096 13342
rect 3124 13314 3148 13342
rect 3176 13314 3187 13342
rect 2877 12558 3187 13314
rect 2877 12530 2888 12558
rect 2916 12530 2940 12558
rect 2968 12530 2992 12558
rect 3020 12530 3044 12558
rect 3072 12530 3096 12558
rect 3124 12530 3148 12558
rect 3176 12530 3187 12558
rect 2877 11774 3187 12530
rect 2877 11746 2888 11774
rect 2916 11746 2940 11774
rect 2968 11746 2992 11774
rect 3020 11746 3044 11774
rect 3072 11746 3096 11774
rect 3124 11746 3148 11774
rect 3176 11746 3187 11774
rect 2877 10990 3187 11746
rect 2877 10962 2888 10990
rect 2916 10962 2940 10990
rect 2968 10962 2992 10990
rect 3020 10962 3044 10990
rect 3072 10962 3096 10990
rect 3124 10962 3148 10990
rect 3176 10962 3187 10990
rect 2877 10206 3187 10962
rect 2877 10178 2888 10206
rect 2916 10178 2940 10206
rect 2968 10178 2992 10206
rect 3020 10178 3044 10206
rect 3072 10178 3096 10206
rect 3124 10178 3148 10206
rect 3176 10178 3187 10206
rect 2877 9422 3187 10178
rect 2877 9394 2888 9422
rect 2916 9394 2940 9422
rect 2968 9394 2992 9422
rect 3020 9394 3044 9422
rect 3072 9394 3096 9422
rect 3124 9394 3148 9422
rect 3176 9394 3187 9422
rect 2877 8638 3187 9394
rect 2877 8610 2888 8638
rect 2916 8610 2940 8638
rect 2968 8610 2992 8638
rect 3020 8610 3044 8638
rect 3072 8610 3096 8638
rect 3124 8610 3148 8638
rect 3176 8610 3187 8638
rect 2877 7854 3187 8610
rect 2877 7826 2888 7854
rect 2916 7826 2940 7854
rect 2968 7826 2992 7854
rect 3020 7826 3044 7854
rect 3072 7826 3096 7854
rect 3124 7826 3148 7854
rect 3176 7826 3187 7854
rect 2877 7070 3187 7826
rect 2877 7042 2888 7070
rect 2916 7042 2940 7070
rect 2968 7042 2992 7070
rect 3020 7042 3044 7070
rect 3072 7042 3096 7070
rect 3124 7042 3148 7070
rect 3176 7042 3187 7070
rect 2877 6286 3187 7042
rect 2877 6258 2888 6286
rect 2916 6258 2940 6286
rect 2968 6258 2992 6286
rect 3020 6258 3044 6286
rect 3072 6258 3096 6286
rect 3124 6258 3148 6286
rect 3176 6258 3187 6286
rect 2877 5502 3187 6258
rect 2877 5474 2888 5502
rect 2916 5474 2940 5502
rect 2968 5474 2992 5502
rect 3020 5474 3044 5502
rect 3072 5474 3096 5502
rect 3124 5474 3148 5502
rect 3176 5474 3187 5502
rect 2877 4718 3187 5474
rect 2877 4690 2888 4718
rect 2916 4690 2940 4718
rect 2968 4690 2992 4718
rect 3020 4690 3044 4718
rect 3072 4690 3096 4718
rect 3124 4690 3148 4718
rect 3176 4690 3187 4718
rect 2877 3934 3187 4690
rect 2877 3906 2888 3934
rect 2916 3906 2940 3934
rect 2968 3906 2992 3934
rect 3020 3906 3044 3934
rect 3072 3906 3096 3934
rect 3124 3906 3148 3934
rect 3176 3906 3187 3934
rect 2877 3150 3187 3906
rect 2877 3122 2888 3150
rect 2916 3122 2940 3150
rect 2968 3122 2992 3150
rect 3020 3122 3044 3150
rect 3072 3122 3096 3150
rect 3124 3122 3148 3150
rect 3176 3122 3187 3150
rect 2877 2366 3187 3122
rect 2877 2338 2888 2366
rect 2916 2338 2940 2366
rect 2968 2338 2992 2366
rect 3020 2338 3044 2366
rect 3072 2338 3096 2366
rect 3124 2338 3148 2366
rect 3176 2338 3187 2366
rect 2877 1582 3187 2338
rect 2877 1554 2888 1582
rect 2916 1554 2940 1582
rect 2968 1554 2992 1582
rect 3020 1554 3044 1582
rect 3072 1554 3096 1582
rect 3124 1554 3148 1582
rect 3176 1554 3187 1582
rect 2877 1538 3187 1554
rect 19017 23142 19327 23158
rect 19017 23114 19028 23142
rect 19056 23114 19080 23142
rect 19108 23114 19132 23142
rect 19160 23114 19184 23142
rect 19212 23114 19236 23142
rect 19264 23114 19288 23142
rect 19316 23114 19327 23142
rect 19017 22358 19327 23114
rect 19017 22330 19028 22358
rect 19056 22330 19080 22358
rect 19108 22330 19132 22358
rect 19160 22330 19184 22358
rect 19212 22330 19236 22358
rect 19264 22330 19288 22358
rect 19316 22330 19327 22358
rect 19017 21574 19327 22330
rect 19017 21546 19028 21574
rect 19056 21546 19080 21574
rect 19108 21546 19132 21574
rect 19160 21546 19184 21574
rect 19212 21546 19236 21574
rect 19264 21546 19288 21574
rect 19316 21546 19327 21574
rect 19017 20790 19327 21546
rect 19017 20762 19028 20790
rect 19056 20762 19080 20790
rect 19108 20762 19132 20790
rect 19160 20762 19184 20790
rect 19212 20762 19236 20790
rect 19264 20762 19288 20790
rect 19316 20762 19327 20790
rect 19017 20006 19327 20762
rect 19017 19978 19028 20006
rect 19056 19978 19080 20006
rect 19108 19978 19132 20006
rect 19160 19978 19184 20006
rect 19212 19978 19236 20006
rect 19264 19978 19288 20006
rect 19316 19978 19327 20006
rect 19017 19222 19327 19978
rect 19017 19194 19028 19222
rect 19056 19194 19080 19222
rect 19108 19194 19132 19222
rect 19160 19194 19184 19222
rect 19212 19194 19236 19222
rect 19264 19194 19288 19222
rect 19316 19194 19327 19222
rect 19017 18438 19327 19194
rect 19017 18410 19028 18438
rect 19056 18410 19080 18438
rect 19108 18410 19132 18438
rect 19160 18410 19184 18438
rect 19212 18410 19236 18438
rect 19264 18410 19288 18438
rect 19316 18410 19327 18438
rect 19017 17654 19327 18410
rect 19017 17626 19028 17654
rect 19056 17626 19080 17654
rect 19108 17626 19132 17654
rect 19160 17626 19184 17654
rect 19212 17626 19236 17654
rect 19264 17626 19288 17654
rect 19316 17626 19327 17654
rect 19017 16870 19327 17626
rect 19017 16842 19028 16870
rect 19056 16842 19080 16870
rect 19108 16842 19132 16870
rect 19160 16842 19184 16870
rect 19212 16842 19236 16870
rect 19264 16842 19288 16870
rect 19316 16842 19327 16870
rect 19017 16086 19327 16842
rect 19017 16058 19028 16086
rect 19056 16058 19080 16086
rect 19108 16058 19132 16086
rect 19160 16058 19184 16086
rect 19212 16058 19236 16086
rect 19264 16058 19288 16086
rect 19316 16058 19327 16086
rect 19017 15302 19327 16058
rect 19017 15274 19028 15302
rect 19056 15274 19080 15302
rect 19108 15274 19132 15302
rect 19160 15274 19184 15302
rect 19212 15274 19236 15302
rect 19264 15274 19288 15302
rect 19316 15274 19327 15302
rect 19017 14518 19327 15274
rect 19017 14490 19028 14518
rect 19056 14490 19080 14518
rect 19108 14490 19132 14518
rect 19160 14490 19184 14518
rect 19212 14490 19236 14518
rect 19264 14490 19288 14518
rect 19316 14490 19327 14518
rect 19017 13734 19327 14490
rect 19017 13706 19028 13734
rect 19056 13706 19080 13734
rect 19108 13706 19132 13734
rect 19160 13706 19184 13734
rect 19212 13706 19236 13734
rect 19264 13706 19288 13734
rect 19316 13706 19327 13734
rect 19017 12950 19327 13706
rect 19017 12922 19028 12950
rect 19056 12922 19080 12950
rect 19108 12922 19132 12950
rect 19160 12922 19184 12950
rect 19212 12922 19236 12950
rect 19264 12922 19288 12950
rect 19316 12922 19327 12950
rect 19017 12166 19327 12922
rect 19017 12138 19028 12166
rect 19056 12138 19080 12166
rect 19108 12138 19132 12166
rect 19160 12138 19184 12166
rect 19212 12138 19236 12166
rect 19264 12138 19288 12166
rect 19316 12138 19327 12166
rect 19017 11382 19327 12138
rect 19017 11354 19028 11382
rect 19056 11354 19080 11382
rect 19108 11354 19132 11382
rect 19160 11354 19184 11382
rect 19212 11354 19236 11382
rect 19264 11354 19288 11382
rect 19316 11354 19327 11382
rect 19017 10598 19327 11354
rect 19017 10570 19028 10598
rect 19056 10570 19080 10598
rect 19108 10570 19132 10598
rect 19160 10570 19184 10598
rect 19212 10570 19236 10598
rect 19264 10570 19288 10598
rect 19316 10570 19327 10598
rect 19017 9814 19327 10570
rect 19017 9786 19028 9814
rect 19056 9786 19080 9814
rect 19108 9786 19132 9814
rect 19160 9786 19184 9814
rect 19212 9786 19236 9814
rect 19264 9786 19288 9814
rect 19316 9786 19327 9814
rect 19017 9030 19327 9786
rect 19017 9002 19028 9030
rect 19056 9002 19080 9030
rect 19108 9002 19132 9030
rect 19160 9002 19184 9030
rect 19212 9002 19236 9030
rect 19264 9002 19288 9030
rect 19316 9002 19327 9030
rect 19017 8246 19327 9002
rect 19017 8218 19028 8246
rect 19056 8218 19080 8246
rect 19108 8218 19132 8246
rect 19160 8218 19184 8246
rect 19212 8218 19236 8246
rect 19264 8218 19288 8246
rect 19316 8218 19327 8246
rect 19017 7462 19327 8218
rect 19017 7434 19028 7462
rect 19056 7434 19080 7462
rect 19108 7434 19132 7462
rect 19160 7434 19184 7462
rect 19212 7434 19236 7462
rect 19264 7434 19288 7462
rect 19316 7434 19327 7462
rect 19017 6678 19327 7434
rect 19017 6650 19028 6678
rect 19056 6650 19080 6678
rect 19108 6650 19132 6678
rect 19160 6650 19184 6678
rect 19212 6650 19236 6678
rect 19264 6650 19288 6678
rect 19316 6650 19327 6678
rect 19017 5894 19327 6650
rect 19017 5866 19028 5894
rect 19056 5866 19080 5894
rect 19108 5866 19132 5894
rect 19160 5866 19184 5894
rect 19212 5866 19236 5894
rect 19264 5866 19288 5894
rect 19316 5866 19327 5894
rect 19017 5110 19327 5866
rect 19017 5082 19028 5110
rect 19056 5082 19080 5110
rect 19108 5082 19132 5110
rect 19160 5082 19184 5110
rect 19212 5082 19236 5110
rect 19264 5082 19288 5110
rect 19316 5082 19327 5110
rect 19017 4326 19327 5082
rect 19017 4298 19028 4326
rect 19056 4298 19080 4326
rect 19108 4298 19132 4326
rect 19160 4298 19184 4326
rect 19212 4298 19236 4326
rect 19264 4298 19288 4326
rect 19316 4298 19327 4326
rect 19017 3542 19327 4298
rect 19017 3514 19028 3542
rect 19056 3514 19080 3542
rect 19108 3514 19132 3542
rect 19160 3514 19184 3542
rect 19212 3514 19236 3542
rect 19264 3514 19288 3542
rect 19316 3514 19327 3542
rect 19017 2758 19327 3514
rect 19017 2730 19028 2758
rect 19056 2730 19080 2758
rect 19108 2730 19132 2758
rect 19160 2730 19184 2758
rect 19212 2730 19236 2758
rect 19264 2730 19288 2758
rect 19316 2730 19327 2758
rect 19017 1974 19327 2730
rect 19017 1946 19028 1974
rect 19056 1946 19080 1974
rect 19108 1946 19132 1974
rect 19160 1946 19184 1974
rect 19212 1946 19236 1974
rect 19264 1946 19288 1974
rect 19316 1946 19327 1974
rect 19017 1538 19327 1946
rect 20877 22750 21187 23158
rect 20877 22722 20888 22750
rect 20916 22722 20940 22750
rect 20968 22722 20992 22750
rect 21020 22722 21044 22750
rect 21072 22722 21096 22750
rect 21124 22722 21148 22750
rect 21176 22722 21187 22750
rect 20877 21966 21187 22722
rect 20877 21938 20888 21966
rect 20916 21938 20940 21966
rect 20968 21938 20992 21966
rect 21020 21938 21044 21966
rect 21072 21938 21096 21966
rect 21124 21938 21148 21966
rect 21176 21938 21187 21966
rect 20877 21182 21187 21938
rect 20877 21154 20888 21182
rect 20916 21154 20940 21182
rect 20968 21154 20992 21182
rect 21020 21154 21044 21182
rect 21072 21154 21096 21182
rect 21124 21154 21148 21182
rect 21176 21154 21187 21182
rect 20877 20398 21187 21154
rect 20877 20370 20888 20398
rect 20916 20370 20940 20398
rect 20968 20370 20992 20398
rect 21020 20370 21044 20398
rect 21072 20370 21096 20398
rect 21124 20370 21148 20398
rect 21176 20370 21187 20398
rect 20877 19614 21187 20370
rect 20877 19586 20888 19614
rect 20916 19586 20940 19614
rect 20968 19586 20992 19614
rect 21020 19586 21044 19614
rect 21072 19586 21096 19614
rect 21124 19586 21148 19614
rect 21176 19586 21187 19614
rect 20877 18830 21187 19586
rect 20877 18802 20888 18830
rect 20916 18802 20940 18830
rect 20968 18802 20992 18830
rect 21020 18802 21044 18830
rect 21072 18802 21096 18830
rect 21124 18802 21148 18830
rect 21176 18802 21187 18830
rect 20877 18046 21187 18802
rect 20877 18018 20888 18046
rect 20916 18018 20940 18046
rect 20968 18018 20992 18046
rect 21020 18018 21044 18046
rect 21072 18018 21096 18046
rect 21124 18018 21148 18046
rect 21176 18018 21187 18046
rect 20877 17262 21187 18018
rect 20877 17234 20888 17262
rect 20916 17234 20940 17262
rect 20968 17234 20992 17262
rect 21020 17234 21044 17262
rect 21072 17234 21096 17262
rect 21124 17234 21148 17262
rect 21176 17234 21187 17262
rect 20877 16478 21187 17234
rect 20877 16450 20888 16478
rect 20916 16450 20940 16478
rect 20968 16450 20992 16478
rect 21020 16450 21044 16478
rect 21072 16450 21096 16478
rect 21124 16450 21148 16478
rect 21176 16450 21187 16478
rect 20877 15694 21187 16450
rect 20877 15666 20888 15694
rect 20916 15666 20940 15694
rect 20968 15666 20992 15694
rect 21020 15666 21044 15694
rect 21072 15666 21096 15694
rect 21124 15666 21148 15694
rect 21176 15666 21187 15694
rect 20877 14910 21187 15666
rect 20877 14882 20888 14910
rect 20916 14882 20940 14910
rect 20968 14882 20992 14910
rect 21020 14882 21044 14910
rect 21072 14882 21096 14910
rect 21124 14882 21148 14910
rect 21176 14882 21187 14910
rect 20877 14126 21187 14882
rect 20877 14098 20888 14126
rect 20916 14098 20940 14126
rect 20968 14098 20992 14126
rect 21020 14098 21044 14126
rect 21072 14098 21096 14126
rect 21124 14098 21148 14126
rect 21176 14098 21187 14126
rect 20877 13342 21187 14098
rect 20877 13314 20888 13342
rect 20916 13314 20940 13342
rect 20968 13314 20992 13342
rect 21020 13314 21044 13342
rect 21072 13314 21096 13342
rect 21124 13314 21148 13342
rect 21176 13314 21187 13342
rect 20877 12558 21187 13314
rect 20877 12530 20888 12558
rect 20916 12530 20940 12558
rect 20968 12530 20992 12558
rect 21020 12530 21044 12558
rect 21072 12530 21096 12558
rect 21124 12530 21148 12558
rect 21176 12530 21187 12558
rect 20877 11774 21187 12530
rect 20877 11746 20888 11774
rect 20916 11746 20940 11774
rect 20968 11746 20992 11774
rect 21020 11746 21044 11774
rect 21072 11746 21096 11774
rect 21124 11746 21148 11774
rect 21176 11746 21187 11774
rect 20877 10990 21187 11746
rect 20877 10962 20888 10990
rect 20916 10962 20940 10990
rect 20968 10962 20992 10990
rect 21020 10962 21044 10990
rect 21072 10962 21096 10990
rect 21124 10962 21148 10990
rect 21176 10962 21187 10990
rect 20877 10206 21187 10962
rect 20877 10178 20888 10206
rect 20916 10178 20940 10206
rect 20968 10178 20992 10206
rect 21020 10178 21044 10206
rect 21072 10178 21096 10206
rect 21124 10178 21148 10206
rect 21176 10178 21187 10206
rect 20877 9422 21187 10178
rect 20877 9394 20888 9422
rect 20916 9394 20940 9422
rect 20968 9394 20992 9422
rect 21020 9394 21044 9422
rect 21072 9394 21096 9422
rect 21124 9394 21148 9422
rect 21176 9394 21187 9422
rect 20877 8638 21187 9394
rect 20877 8610 20888 8638
rect 20916 8610 20940 8638
rect 20968 8610 20992 8638
rect 21020 8610 21044 8638
rect 21072 8610 21096 8638
rect 21124 8610 21148 8638
rect 21176 8610 21187 8638
rect 20877 7854 21187 8610
rect 20877 7826 20888 7854
rect 20916 7826 20940 7854
rect 20968 7826 20992 7854
rect 21020 7826 21044 7854
rect 21072 7826 21096 7854
rect 21124 7826 21148 7854
rect 21176 7826 21187 7854
rect 20877 7070 21187 7826
rect 20877 7042 20888 7070
rect 20916 7042 20940 7070
rect 20968 7042 20992 7070
rect 21020 7042 21044 7070
rect 21072 7042 21096 7070
rect 21124 7042 21148 7070
rect 21176 7042 21187 7070
rect 20877 6286 21187 7042
rect 20877 6258 20888 6286
rect 20916 6258 20940 6286
rect 20968 6258 20992 6286
rect 21020 6258 21044 6286
rect 21072 6258 21096 6286
rect 21124 6258 21148 6286
rect 21176 6258 21187 6286
rect 20877 5502 21187 6258
rect 20877 5474 20888 5502
rect 20916 5474 20940 5502
rect 20968 5474 20992 5502
rect 21020 5474 21044 5502
rect 21072 5474 21096 5502
rect 21124 5474 21148 5502
rect 21176 5474 21187 5502
rect 20877 4718 21187 5474
rect 20877 4690 20888 4718
rect 20916 4690 20940 4718
rect 20968 4690 20992 4718
rect 21020 4690 21044 4718
rect 21072 4690 21096 4718
rect 21124 4690 21148 4718
rect 21176 4690 21187 4718
rect 20877 3934 21187 4690
rect 20877 3906 20888 3934
rect 20916 3906 20940 3934
rect 20968 3906 20992 3934
rect 21020 3906 21044 3934
rect 21072 3906 21096 3934
rect 21124 3906 21148 3934
rect 21176 3906 21187 3934
rect 20877 3150 21187 3906
rect 20877 3122 20888 3150
rect 20916 3122 20940 3150
rect 20968 3122 20992 3150
rect 21020 3122 21044 3150
rect 21072 3122 21096 3150
rect 21124 3122 21148 3150
rect 21176 3122 21187 3150
rect 20877 2366 21187 3122
rect 20877 2338 20888 2366
rect 20916 2338 20940 2366
rect 20968 2338 20992 2366
rect 21020 2338 21044 2366
rect 21072 2338 21096 2366
rect 21124 2338 21148 2366
rect 21176 2338 21187 2366
rect 20877 1582 21187 2338
rect 20877 1554 20888 1582
rect 20916 1554 20940 1582
rect 20968 1554 20992 1582
rect 21020 1554 21044 1582
rect 21072 1554 21096 1582
rect 21124 1554 21148 1582
rect 21176 1554 21187 1582
rect 20877 1538 21187 1554
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1__I1 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 13272 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3__D
timestamp 1666464484
transform 1 0 13552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_core_clock_I
timestamp 1666464484
transform -1 0 12544 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_0__f_core_clock_I
timestamp 1666464484
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_1__f_core_clock_I
timestamp 1666464484
transform 1 0 16240 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1666464484
transform -1 0 18648 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output2_I
timestamp 1666464484
transform -1 0 1400 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 2576 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37
timestamp 1666464484
transform 1 0 2744 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1666464484
transform 1 0 4536 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72
timestamp 1666464484
transform 1 0 4704 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1666464484
transform 1 0 6496 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_107
timestamp 1666464484
transform 1 0 6664 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1666464484
transform 1 0 8456 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_142
timestamp 1666464484
transform 1 0 8624 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1666464484
transform 1 0 10416 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_177
timestamp 1666464484
transform 1 0 10584 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1666464484
transform 1 0 12376 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_212
timestamp 1666464484
transform 1 0 12544 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1666464484
transform 1 0 14336 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_247
timestamp 1666464484
transform 1 0 14504 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1666464484
transform 1 0 16296 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_282
timestamp 1666464484
transform 1 0 16464 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1666464484
transform 1 0 18256 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_317 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 18424 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_321
timestamp 1666464484
transform 1 0 18648 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_329 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 19096 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_345 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 19992 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1666464484
transform 1 0 20216 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_352
timestamp 1666464484
transform 1 0 20384 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1666464484
transform 1 0 22176 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_387
timestamp 1666464484
transform 1 0 22344 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1666464484
transform 1 0 24136 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1666464484
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1666464484
transform 1 0 4592 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_73
timestamp 1666464484
transform 1 0 4760 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_137
timestamp 1666464484
transform 1 0 8344 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1666464484
transform 1 0 8568 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_144
timestamp 1666464484
transform 1 0 8736 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_208
timestamp 1666464484
transform 1 0 12320 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1666464484
transform 1 0 12544 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_215
timestamp 1666464484
transform 1 0 12712 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_279
timestamp 1666464484
transform 1 0 16296 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1666464484
transform 1 0 16520 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_286
timestamp 1666464484
transform 1 0 16688 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_350
timestamp 1666464484
transform 1 0 20272 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1666464484
transform 1 0 20496 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_357
timestamp 1666464484
transform 1 0 20664 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_389
timestamp 1666464484
transform 1 0 22456 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_405 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 23352 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_413
timestamp 1666464484
transform 1 0 23800 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_417
timestamp 1666464484
transform 1 0 24024 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_419
timestamp 1666464484
transform 1 0 24136 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1666464484
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1666464484
transform 1 0 2576 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1666464484
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1666464484
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1666464484
transform 1 0 6552 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108
timestamp 1666464484
transform 1 0 6720 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1666464484
transform 1 0 10304 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1666464484
transform 1 0 10528 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_179
timestamp 1666464484
transform 1 0 10696 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_243
timestamp 1666464484
transform 1 0 14280 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1666464484
transform 1 0 14504 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_250
timestamp 1666464484
transform 1 0 14672 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_314
timestamp 1666464484
transform 1 0 18256 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1666464484
transform 1 0 18480 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_321
timestamp 1666464484
transform 1 0 18648 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_385
timestamp 1666464484
transform 1 0 22232 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1666464484
transform 1 0 22456 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_392
timestamp 1666464484
transform 1 0 22624 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_408
timestamp 1666464484
transform 1 0 23520 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_416
timestamp 1666464484
transform 1 0 23968 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1666464484
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1666464484
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1666464484
transform 1 0 4592 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1666464484
transform 1 0 4760 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1666464484
transform 1 0 8344 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1666464484
transform 1 0 8568 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1666464484
transform 1 0 8736 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1666464484
transform 1 0 12320 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1666464484
transform 1 0 12544 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1666464484
transform 1 0 12712 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1666464484
transform 1 0 16296 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1666464484
transform 1 0 16520 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1666464484
transform 1 0 16688 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_350
timestamp 1666464484
transform 1 0 20272 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1666464484
transform 1 0 20496 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_357
timestamp 1666464484
transform 1 0 20664 0 -1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_389
timestamp 1666464484
transform 1 0 22456 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_405
timestamp 1666464484
transform 1 0 23352 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_413
timestamp 1666464484
transform 1 0 23800 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_417
timestamp 1666464484
transform 1 0 24024 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_419
timestamp 1666464484
transform 1 0 24136 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1666464484
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1666464484
transform 1 0 2576 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1666464484
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1666464484
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1666464484
transform 1 0 6552 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1666464484
transform 1 0 6720 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1666464484
transform 1 0 10304 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1666464484
transform 1 0 10528 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1666464484
transform 1 0 10696 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1666464484
transform 1 0 14280 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1666464484
transform 1 0 14504 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1666464484
transform 1 0 14672 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1666464484
transform 1 0 18256 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1666464484
transform 1 0 18480 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1666464484
transform 1 0 18648 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1666464484
transform 1 0 22232 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1666464484
transform 1 0 22456 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_392
timestamp 1666464484
transform 1 0 22624 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_408
timestamp 1666464484
transform 1 0 23520 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_416
timestamp 1666464484
transform 1 0 23968 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1666464484
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1666464484
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1666464484
transform 1 0 4592 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1666464484
transform 1 0 4760 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1666464484
transform 1 0 8344 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1666464484
transform 1 0 8568 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_144
timestamp 1666464484
transform 1 0 8736 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_152
timestamp 1666464484
transform 1 0 9184 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_156
timestamp 1666464484
transform 1 0 9408 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_208
timestamp 1666464484
transform 1 0 12320 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1666464484
transform 1 0 12544 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1666464484
transform 1 0 12712 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1666464484
transform 1 0 16296 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1666464484
transform 1 0 16520 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1666464484
transform 1 0 16688 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1666464484
transform 1 0 20272 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1666464484
transform 1 0 20496 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_357
timestamp 1666464484
transform 1 0 20664 0 -1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_389
timestamp 1666464484
transform 1 0 22456 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_405
timestamp 1666464484
transform 1 0 23352 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_413
timestamp 1666464484
transform 1 0 23800 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_417
timestamp 1666464484
transform 1 0 24024 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_419
timestamp 1666464484
transform 1 0 24136 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1666464484
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1666464484
transform 1 0 2576 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1666464484
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1666464484
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1666464484
transform 1 0 6552 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1666464484
transform 1 0 6720 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1666464484
transform 1 0 10304 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1666464484
transform 1 0 10528 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1666464484
transform 1 0 10696 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1666464484
transform 1 0 14280 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1666464484
transform 1 0 14504 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1666464484
transform 1 0 14672 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1666464484
transform 1 0 18256 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1666464484
transform 1 0 18480 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1666464484
transform 1 0 18648 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1666464484
transform 1 0 22232 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1666464484
transform 1 0 22456 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_392
timestamp 1666464484
transform 1 0 22624 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_408
timestamp 1666464484
transform 1 0 23520 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_416
timestamp 1666464484
transform 1 0 23968 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_2
timestamp 1666464484
transform 1 0 784 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_9
timestamp 1666464484
transform 1 0 1176 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_13
timestamp 1666464484
transform 1 0 1400 0 -1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_45
timestamp 1666464484
transform 1 0 3192 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_61
timestamp 1666464484
transform 1 0 4088 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_69
timestamp 1666464484
transform 1 0 4536 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1666464484
transform 1 0 4760 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1666464484
transform 1 0 8344 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1666464484
transform 1 0 8568 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1666464484
transform 1 0 8736 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1666464484
transform 1 0 12320 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1666464484
transform 1 0 12544 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1666464484
transform 1 0 12712 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1666464484
transform 1 0 16296 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1666464484
transform 1 0 16520 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1666464484
transform 1 0 16688 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1666464484
transform 1 0 20272 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1666464484
transform 1 0 20496 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_357
timestamp 1666464484
transform 1 0 20664 0 -1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_389
timestamp 1666464484
transform 1 0 22456 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_405
timestamp 1666464484
transform 1 0 23352 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_413
timestamp 1666464484
transform 1 0 23800 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_417
timestamp 1666464484
transform 1 0 24024 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_419
timestamp 1666464484
transform 1 0 24136 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1666464484
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1666464484
transform 1 0 2576 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1666464484
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1666464484
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1666464484
transform 1 0 6552 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1666464484
transform 1 0 6720 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1666464484
transform 1 0 10304 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1666464484
transform 1 0 10528 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_179
timestamp 1666464484
transform 1 0 10696 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_195
timestamp 1666464484
transform 1 0 11592 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_228
timestamp 1666464484
transform 1 0 13440 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_232
timestamp 1666464484
transform 1 0 13664 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1666464484
transform 1 0 14672 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1666464484
transform 1 0 18256 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1666464484
transform 1 0 18480 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1666464484
transform 1 0 18648 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1666464484
transform 1 0 22232 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1666464484
transform 1 0 22456 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_392
timestamp 1666464484
transform 1 0 22624 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_408
timestamp 1666464484
transform 1 0 23520 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_416
timestamp 1666464484
transform 1 0 23968 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1666464484
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1666464484
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1666464484
transform 1 0 4592 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1666464484
transform 1 0 4760 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1666464484
transform 1 0 8344 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1666464484
transform 1 0 8568 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_144
timestamp 1666464484
transform 1 0 8736 0 -1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_176
timestamp 1666464484
transform 1 0 10528 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_192
timestamp 1666464484
transform 1 0 11424 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_202
timestamp 1666464484
transform 1 0 11984 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1666464484
transform 1 0 12544 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_215
timestamp 1666464484
transform 1 0 12712 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_266
timestamp 1666464484
transform 1 0 15568 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_282
timestamp 1666464484
transform 1 0 16464 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1666464484
transform 1 0 16688 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1666464484
transform 1 0 20272 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1666464484
transform 1 0 20496 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_357
timestamp 1666464484
transform 1 0 20664 0 -1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_389
timestamp 1666464484
transform 1 0 22456 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_405
timestamp 1666464484
transform 1 0 23352 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_413
timestamp 1666464484
transform 1 0 23800 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_417
timestamp 1666464484
transform 1 0 24024 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_419
timestamp 1666464484
transform 1 0 24136 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1666464484
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1666464484
transform 1 0 2576 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1666464484
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1666464484
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1666464484
transform 1 0 6552 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1666464484
transform 1 0 6720 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1666464484
transform 1 0 10304 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1666464484
transform 1 0 10528 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_179
timestamp 1666464484
transform 1 0 10696 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_195
timestamp 1666464484
transform 1 0 11592 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_203
timestamp 1666464484
transform 1 0 12040 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_205
timestamp 1666464484
transform 1 0 12152 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_221
timestamp 1666464484
transform 1 0 13048 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_225
timestamp 1666464484
transform 1 0 13272 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_241
timestamp 1666464484
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_245
timestamp 1666464484
transform 1 0 14392 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1666464484
transform 1 0 14504 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1666464484
transform 1 0 14672 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1666464484
transform 1 0 18256 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1666464484
transform 1 0 18480 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1666464484
transform 1 0 18648 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1666464484
transform 1 0 22232 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1666464484
transform 1 0 22456 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_392
timestamp 1666464484
transform 1 0 22624 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_408
timestamp 1666464484
transform 1 0 23520 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_416
timestamp 1666464484
transform 1 0 23968 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1666464484
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1666464484
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1666464484
transform 1 0 4592 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1666464484
transform 1 0 4760 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1666464484
transform 1 0 8344 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1666464484
transform 1 0 8568 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1666464484
transform 1 0 8736 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1666464484
transform 1 0 12320 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1666464484
transform 1 0 12544 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_215
timestamp 1666464484
transform 1 0 12712 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_223
timestamp 1666464484
transform 1 0 13160 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_225
timestamp 1666464484
transform 1 0 13272 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_276
timestamp 1666464484
transform 1 0 16128 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_280
timestamp 1666464484
transform 1 0 16352 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1666464484
transform 1 0 16688 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1666464484
transform 1 0 20272 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1666464484
transform 1 0 20496 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_357
timestamp 1666464484
transform 1 0 20664 0 -1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_389
timestamp 1666464484
transform 1 0 22456 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_405
timestamp 1666464484
transform 1 0 23352 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_413
timestamp 1666464484
transform 1 0 23800 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_417
timestamp 1666464484
transform 1 0 24024 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_419
timestamp 1666464484
transform 1 0 24136 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1666464484
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1666464484
transform 1 0 2576 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1666464484
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1666464484
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1666464484
transform 1 0 6552 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1666464484
transform 1 0 6720 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1666464484
transform 1 0 10304 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1666464484
transform 1 0 10528 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1666464484
transform 1 0 10696 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1666464484
transform 1 0 14280 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1666464484
transform 1 0 14504 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1666464484
transform 1 0 14672 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1666464484
transform 1 0 18256 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1666464484
transform 1 0 18480 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1666464484
transform 1 0 18648 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1666464484
transform 1 0 22232 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1666464484
transform 1 0 22456 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_392
timestamp 1666464484
transform 1 0 22624 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_408
timestamp 1666464484
transform 1 0 23520 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_416
timestamp 1666464484
transform 1 0 23968 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1666464484
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1666464484
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1666464484
transform 1 0 4592 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1666464484
transform 1 0 4760 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1666464484
transform 1 0 8344 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1666464484
transform 1 0 8568 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1666464484
transform 1 0 8736 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1666464484
transform 1 0 12320 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1666464484
transform 1 0 12544 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1666464484
transform 1 0 12712 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1666464484
transform 1 0 16296 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1666464484
transform 1 0 16520 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1666464484
transform 1 0 16688 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1666464484
transform 1 0 20272 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1666464484
transform 1 0 20496 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_357
timestamp 1666464484
transform 1 0 20664 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_389
timestamp 1666464484
transform 1 0 22456 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_405
timestamp 1666464484
transform 1 0 23352 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_413
timestamp 1666464484
transform 1 0 23800 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_417
timestamp 1666464484
transform 1 0 24024 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_419
timestamp 1666464484
transform 1 0 24136 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1666464484
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1666464484
transform 1 0 2576 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1666464484
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1666464484
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1666464484
transform 1 0 6552 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1666464484
transform 1 0 6720 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1666464484
transform 1 0 10304 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1666464484
transform 1 0 10528 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1666464484
transform 1 0 10696 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1666464484
transform 1 0 14280 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1666464484
transform 1 0 14504 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1666464484
transform 1 0 14672 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1666464484
transform 1 0 18256 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1666464484
transform 1 0 18480 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1666464484
transform 1 0 18648 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1666464484
transform 1 0 22232 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1666464484
transform 1 0 22456 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_392
timestamp 1666464484
transform 1 0 22624 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_408
timestamp 1666464484
transform 1 0 23520 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_416
timestamp 1666464484
transform 1 0 23968 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1666464484
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1666464484
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1666464484
transform 1 0 4592 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1666464484
transform 1 0 4760 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1666464484
transform 1 0 8344 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1666464484
transform 1 0 8568 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1666464484
transform 1 0 8736 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1666464484
transform 1 0 12320 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1666464484
transform 1 0 12544 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1666464484
transform 1 0 12712 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1666464484
transform 1 0 16296 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1666464484
transform 1 0 16520 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1666464484
transform 1 0 16688 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1666464484
transform 1 0 20272 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1666464484
transform 1 0 20496 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_357
timestamp 1666464484
transform 1 0 20664 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_389
timestamp 1666464484
transform 1 0 22456 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_405
timestamp 1666464484
transform 1 0 23352 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_413
timestamp 1666464484
transform 1 0 23800 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_417
timestamp 1666464484
transform 1 0 24024 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_419
timestamp 1666464484
transform 1 0 24136 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1666464484
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1666464484
transform 1 0 2576 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1666464484
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1666464484
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1666464484
transform 1 0 6552 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1666464484
transform 1 0 6720 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1666464484
transform 1 0 10304 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1666464484
transform 1 0 10528 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1666464484
transform 1 0 10696 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1666464484
transform 1 0 14280 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1666464484
transform 1 0 14504 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1666464484
transform 1 0 14672 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1666464484
transform 1 0 18256 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1666464484
transform 1 0 18480 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1666464484
transform 1 0 18648 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1666464484
transform 1 0 22232 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1666464484
transform 1 0 22456 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_392
timestamp 1666464484
transform 1 0 22624 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_408
timestamp 1666464484
transform 1 0 23520 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_416
timestamp 1666464484
transform 1 0 23968 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1666464484
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1666464484
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1666464484
transform 1 0 4592 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1666464484
transform 1 0 4760 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1666464484
transform 1 0 8344 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1666464484
transform 1 0 8568 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1666464484
transform 1 0 8736 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1666464484
transform 1 0 12320 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1666464484
transform 1 0 12544 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1666464484
transform 1 0 12712 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1666464484
transform 1 0 16296 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1666464484
transform 1 0 16520 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1666464484
transform 1 0 16688 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1666464484
transform 1 0 20272 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1666464484
transform 1 0 20496 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_357
timestamp 1666464484
transform 1 0 20664 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_389
timestamp 1666464484
transform 1 0 22456 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_405
timestamp 1666464484
transform 1 0 23352 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_413
timestamp 1666464484
transform 1 0 23800 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_417
timestamp 1666464484
transform 1 0 24024 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_419
timestamp 1666464484
transform 1 0 24136 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_2
timestamp 1666464484
transform 1 0 784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1666464484
transform 1 0 2576 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1666464484
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1666464484
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1666464484
transform 1 0 6552 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1666464484
transform 1 0 6720 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1666464484
transform 1 0 10304 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1666464484
transform 1 0 10528 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1666464484
transform 1 0 10696 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1666464484
transform 1 0 14280 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1666464484
transform 1 0 14504 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1666464484
transform 1 0 14672 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1666464484
transform 1 0 18256 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1666464484
transform 1 0 18480 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1666464484
transform 1 0 18648 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1666464484
transform 1 0 22232 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1666464484
transform 1 0 22456 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_392
timestamp 1666464484
transform 1 0 22624 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_408
timestamp 1666464484
transform 1 0 23520 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_416
timestamp 1666464484
transform 1 0 23968 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1666464484
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1666464484
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1666464484
transform 1 0 4592 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1666464484
transform 1 0 4760 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1666464484
transform 1 0 8344 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1666464484
transform 1 0 8568 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1666464484
transform 1 0 8736 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1666464484
transform 1 0 12320 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1666464484
transform 1 0 12544 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1666464484
transform 1 0 12712 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1666464484
transform 1 0 16296 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1666464484
transform 1 0 16520 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1666464484
transform 1 0 16688 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1666464484
transform 1 0 20272 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1666464484
transform 1 0 20496 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_357
timestamp 1666464484
transform 1 0 20664 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_389
timestamp 1666464484
transform 1 0 22456 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_405
timestamp 1666464484
transform 1 0 23352 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_413
timestamp 1666464484
transform 1 0 23800 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_417
timestamp 1666464484
transform 1 0 24024 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_419
timestamp 1666464484
transform 1 0 24136 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1666464484
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1666464484
transform 1 0 2576 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1666464484
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1666464484
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1666464484
transform 1 0 6552 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1666464484
transform 1 0 6720 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1666464484
transform 1 0 10304 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1666464484
transform 1 0 10528 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1666464484
transform 1 0 10696 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1666464484
transform 1 0 14280 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1666464484
transform 1 0 14504 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1666464484
transform 1 0 14672 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1666464484
transform 1 0 18256 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1666464484
transform 1 0 18480 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1666464484
transform 1 0 18648 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1666464484
transform 1 0 22232 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1666464484
transform 1 0 22456 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_392
timestamp 1666464484
transform 1 0 22624 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_408
timestamp 1666464484
transform 1 0 23520 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_416
timestamp 1666464484
transform 1 0 23968 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1666464484
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1666464484
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1666464484
transform 1 0 4592 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1666464484
transform 1 0 4760 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1666464484
transform 1 0 8344 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1666464484
transform 1 0 8568 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1666464484
transform 1 0 8736 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1666464484
transform 1 0 12320 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1666464484
transform 1 0 12544 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1666464484
transform 1 0 12712 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1666464484
transform 1 0 16296 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1666464484
transform 1 0 16520 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1666464484
transform 1 0 16688 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1666464484
transform 1 0 20272 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1666464484
transform 1 0 20496 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_357
timestamp 1666464484
transform 1 0 20664 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_389
timestamp 1666464484
transform 1 0 22456 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_405
timestamp 1666464484
transform 1 0 23352 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_413
timestamp 1666464484
transform 1 0 23800 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_417
timestamp 1666464484
transform 1 0 24024 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_419
timestamp 1666464484
transform 1 0 24136 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1666464484
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1666464484
transform 1 0 2576 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1666464484
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1666464484
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1666464484
transform 1 0 6552 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1666464484
transform 1 0 6720 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1666464484
transform 1 0 10304 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1666464484
transform 1 0 10528 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1666464484
transform 1 0 10696 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1666464484
transform 1 0 14280 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1666464484
transform 1 0 14504 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1666464484
transform 1 0 14672 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1666464484
transform 1 0 18256 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1666464484
transform 1 0 18480 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1666464484
transform 1 0 18648 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1666464484
transform 1 0 22232 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1666464484
transform 1 0 22456 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_392
timestamp 1666464484
transform 1 0 22624 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_408
timestamp 1666464484
transform 1 0 23520 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_416
timestamp 1666464484
transform 1 0 23968 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_2
timestamp 1666464484
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_66
timestamp 1666464484
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1666464484
transform 1 0 4592 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1666464484
transform 1 0 4760 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1666464484
transform 1 0 8344 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1666464484
transform 1 0 8568 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1666464484
transform 1 0 8736 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1666464484
transform 1 0 12320 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1666464484
transform 1 0 12544 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1666464484
transform 1 0 12712 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1666464484
transform 1 0 16296 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1666464484
transform 1 0 16520 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1666464484
transform 1 0 16688 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1666464484
transform 1 0 20272 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1666464484
transform 1 0 20496 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_357
timestamp 1666464484
transform 1 0 20664 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_389
timestamp 1666464484
transform 1 0 22456 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_405
timestamp 1666464484
transform 1 0 23352 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_413
timestamp 1666464484
transform 1 0 23800 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_417
timestamp 1666464484
transform 1 0 24024 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_419
timestamp 1666464484
transform 1 0 24136 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_2
timestamp 1666464484
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1666464484
transform 1 0 2576 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1666464484
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1666464484
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1666464484
transform 1 0 6552 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1666464484
transform 1 0 6720 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1666464484
transform 1 0 10304 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1666464484
transform 1 0 10528 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1666464484
transform 1 0 10696 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1666464484
transform 1 0 14280 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1666464484
transform 1 0 14504 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1666464484
transform 1 0 14672 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1666464484
transform 1 0 18256 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1666464484
transform 1 0 18480 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1666464484
transform 1 0 18648 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1666464484
transform 1 0 22232 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1666464484
transform 1 0 22456 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_392
timestamp 1666464484
transform 1 0 22624 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_408
timestamp 1666464484
transform 1 0 23520 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_416
timestamp 1666464484
transform 1 0 23968 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_2
timestamp 1666464484
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_66
timestamp 1666464484
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1666464484
transform 1 0 4592 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1666464484
transform 1 0 4760 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1666464484
transform 1 0 8344 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1666464484
transform 1 0 8568 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1666464484
transform 1 0 8736 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1666464484
transform 1 0 12320 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1666464484
transform 1 0 12544 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1666464484
transform 1 0 12712 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1666464484
transform 1 0 16296 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1666464484
transform 1 0 16520 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1666464484
transform 1 0 16688 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1666464484
transform 1 0 20272 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1666464484
transform 1 0 20496 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_357
timestamp 1666464484
transform 1 0 20664 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_389
timestamp 1666464484
transform 1 0 22456 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_405
timestamp 1666464484
transform 1 0 23352 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_413
timestamp 1666464484
transform 1 0 23800 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_417
timestamp 1666464484
transform 1 0 24024 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_419
timestamp 1666464484
transform 1 0 24136 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1666464484
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1666464484
transform 1 0 2576 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1666464484
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1666464484
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1666464484
transform 1 0 6552 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1666464484
transform 1 0 6720 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1666464484
transform 1 0 10304 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1666464484
transform 1 0 10528 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1666464484
transform 1 0 10696 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1666464484
transform 1 0 14280 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1666464484
transform 1 0 14504 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1666464484
transform 1 0 14672 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1666464484
transform 1 0 18256 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1666464484
transform 1 0 18480 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1666464484
transform 1 0 18648 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1666464484
transform 1 0 22232 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1666464484
transform 1 0 22456 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_392
timestamp 1666464484
transform 1 0 22624 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_408
timestamp 1666464484
transform 1 0 23520 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_416
timestamp 1666464484
transform 1 0 23968 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1666464484
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1666464484
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1666464484
transform 1 0 4592 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1666464484
transform 1 0 4760 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1666464484
transform 1 0 8344 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1666464484
transform 1 0 8568 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1666464484
transform 1 0 8736 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1666464484
transform 1 0 12320 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1666464484
transform 1 0 12544 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1666464484
transform 1 0 12712 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1666464484
transform 1 0 16296 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1666464484
transform 1 0 16520 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1666464484
transform 1 0 16688 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1666464484
transform 1 0 20272 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1666464484
transform 1 0 20496 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_357
timestamp 1666464484
transform 1 0 20664 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_389
timestamp 1666464484
transform 1 0 22456 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_405
timestamp 1666464484
transform 1 0 23352 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_413
timestamp 1666464484
transform 1 0 23800 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_417
timestamp 1666464484
transform 1 0 24024 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_419
timestamp 1666464484
transform 1 0 24136 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_2
timestamp 1666464484
transform 1 0 784 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_7
timestamp 1666464484
transform 1 0 1064 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_23
timestamp 1666464484
transform 1 0 1960 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_31
timestamp 1666464484
transform 1 0 2408 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1666464484
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1666464484
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1666464484
transform 1 0 6552 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1666464484
transform 1 0 6720 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1666464484
transform 1 0 10304 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1666464484
transform 1 0 10528 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1666464484
transform 1 0 10696 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1666464484
transform 1 0 14280 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1666464484
transform 1 0 14504 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1666464484
transform 1 0 14672 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1666464484
transform 1 0 18256 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1666464484
transform 1 0 18480 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1666464484
transform 1 0 18648 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1666464484
transform 1 0 22232 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1666464484
transform 1 0 22456 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_392
timestamp 1666464484
transform 1 0 22624 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_408
timestamp 1666464484
transform 1 0 23520 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_416
timestamp 1666464484
transform 1 0 23968 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1666464484
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1666464484
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1666464484
transform 1 0 4592 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1666464484
transform 1 0 4760 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1666464484
transform 1 0 8344 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1666464484
transform 1 0 8568 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1666464484
transform 1 0 8736 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1666464484
transform 1 0 12320 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1666464484
transform 1 0 12544 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1666464484
transform 1 0 12712 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1666464484
transform 1 0 16296 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1666464484
transform 1 0 16520 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1666464484
transform 1 0 16688 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1666464484
transform 1 0 20272 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1666464484
transform 1 0 20496 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_357
timestamp 1666464484
transform 1 0 20664 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_389
timestamp 1666464484
transform 1 0 22456 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_405
timestamp 1666464484
transform 1 0 23352 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_413
timestamp 1666464484
transform 1 0 23800 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_417
timestamp 1666464484
transform 1 0 24024 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_419
timestamp 1666464484
transform 1 0 24136 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1666464484
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1666464484
transform 1 0 2576 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1666464484
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1666464484
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1666464484
transform 1 0 6552 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1666464484
transform 1 0 6720 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1666464484
transform 1 0 10304 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1666464484
transform 1 0 10528 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1666464484
transform 1 0 10696 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1666464484
transform 1 0 14280 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1666464484
transform 1 0 14504 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1666464484
transform 1 0 14672 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1666464484
transform 1 0 18256 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1666464484
transform 1 0 18480 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1666464484
transform 1 0 18648 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1666464484
transform 1 0 22232 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1666464484
transform 1 0 22456 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_392
timestamp 1666464484
transform 1 0 22624 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_408
timestamp 1666464484
transform 1 0 23520 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_416
timestamp 1666464484
transform 1 0 23968 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1666464484
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1666464484
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1666464484
transform 1 0 4592 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1666464484
transform 1 0 4760 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1666464484
transform 1 0 8344 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1666464484
transform 1 0 8568 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1666464484
transform 1 0 8736 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1666464484
transform 1 0 12320 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1666464484
transform 1 0 12544 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1666464484
transform 1 0 12712 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1666464484
transform 1 0 16296 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1666464484
transform 1 0 16520 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1666464484
transform 1 0 16688 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1666464484
transform 1 0 20272 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1666464484
transform 1 0 20496 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_357
timestamp 1666464484
transform 1 0 20664 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_389
timestamp 1666464484
transform 1 0 22456 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_405
timestamp 1666464484
transform 1 0 23352 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_413
timestamp 1666464484
transform 1 0 23800 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_417
timestamp 1666464484
transform 1 0 24024 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_419
timestamp 1666464484
transform 1 0 24136 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_2
timestamp 1666464484
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1666464484
transform 1 0 2576 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1666464484
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1666464484
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1666464484
transform 1 0 6552 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1666464484
transform 1 0 6720 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1666464484
transform 1 0 10304 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1666464484
transform 1 0 10528 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1666464484
transform 1 0 10696 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1666464484
transform 1 0 14280 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1666464484
transform 1 0 14504 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1666464484
transform 1 0 14672 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1666464484
transform 1 0 18256 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1666464484
transform 1 0 18480 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1666464484
transform 1 0 18648 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1666464484
transform 1 0 22232 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1666464484
transform 1 0 22456 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_392
timestamp 1666464484
transform 1 0 22624 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_408
timestamp 1666464484
transform 1 0 23520 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_416
timestamp 1666464484
transform 1 0 23968 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1666464484
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1666464484
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1666464484
transform 1 0 4592 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1666464484
transform 1 0 4760 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1666464484
transform 1 0 8344 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1666464484
transform 1 0 8568 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1666464484
transform 1 0 8736 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1666464484
transform 1 0 12320 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1666464484
transform 1 0 12544 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1666464484
transform 1 0 12712 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1666464484
transform 1 0 16296 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1666464484
transform 1 0 16520 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1666464484
transform 1 0 16688 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1666464484
transform 1 0 20272 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1666464484
transform 1 0 20496 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_357
timestamp 1666464484
transform 1 0 20664 0 -1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_389
timestamp 1666464484
transform 1 0 22456 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_405
timestamp 1666464484
transform 1 0 23352 0 -1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_413
timestamp 1666464484
transform 1 0 23800 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_417
timestamp 1666464484
transform 1 0 24024 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_419
timestamp 1666464484
transform 1 0 24136 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_2
timestamp 1666464484
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1666464484
transform 1 0 2576 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1666464484
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1666464484
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1666464484
transform 1 0 6552 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1666464484
transform 1 0 6720 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1666464484
transform 1 0 10304 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1666464484
transform 1 0 10528 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1666464484
transform 1 0 10696 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1666464484
transform 1 0 14280 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1666464484
transform 1 0 14504 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1666464484
transform 1 0 14672 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1666464484
transform 1 0 18256 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1666464484
transform 1 0 18480 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1666464484
transform 1 0 18648 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1666464484
transform 1 0 22232 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1666464484
transform 1 0 22456 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_392
timestamp 1666464484
transform 1 0 22624 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_408
timestamp 1666464484
transform 1 0 23520 0 1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_416
timestamp 1666464484
transform 1 0 23968 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1666464484
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1666464484
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1666464484
transform 1 0 4592 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1666464484
transform 1 0 4760 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1666464484
transform 1 0 8344 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1666464484
transform 1 0 8568 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1666464484
transform 1 0 8736 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1666464484
transform 1 0 12320 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1666464484
transform 1 0 12544 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1666464484
transform 1 0 12712 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1666464484
transform 1 0 16296 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1666464484
transform 1 0 16520 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1666464484
transform 1 0 16688 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1666464484
transform 1 0 20272 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1666464484
transform 1 0 20496 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_357
timestamp 1666464484
transform 1 0 20664 0 -1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_389
timestamp 1666464484
transform 1 0 22456 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_405
timestamp 1666464484
transform 1 0 23352 0 -1 15680
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_413
timestamp 1666464484
transform 1 0 23800 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_417
timestamp 1666464484
transform 1 0 24024 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_419
timestamp 1666464484
transform 1 0 24136 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1666464484
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1666464484
transform 1 0 2576 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1666464484
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1666464484
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1666464484
transform 1 0 6552 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1666464484
transform 1 0 6720 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1666464484
transform 1 0 10304 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1666464484
transform 1 0 10528 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1666464484
transform 1 0 10696 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1666464484
transform 1 0 14280 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1666464484
transform 1 0 14504 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1666464484
transform 1 0 14672 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1666464484
transform 1 0 18256 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1666464484
transform 1 0 18480 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1666464484
transform 1 0 18648 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1666464484
transform 1 0 22232 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1666464484
transform 1 0 22456 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_392
timestamp 1666464484
transform 1 0 22624 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_408
timestamp 1666464484
transform 1 0 23520 0 1 15680
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_416
timestamp 1666464484
transform 1 0 23968 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1666464484
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1666464484
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1666464484
transform 1 0 4592 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1666464484
transform 1 0 4760 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1666464484
transform 1 0 8344 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1666464484
transform 1 0 8568 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1666464484
transform 1 0 8736 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1666464484
transform 1 0 12320 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1666464484
transform 1 0 12544 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1666464484
transform 1 0 12712 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1666464484
transform 1 0 16296 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1666464484
transform 1 0 16520 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1666464484
transform 1 0 16688 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1666464484
transform 1 0 20272 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1666464484
transform 1 0 20496 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_357
timestamp 1666464484
transform 1 0 20664 0 -1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_389
timestamp 1666464484
transform 1 0 22456 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_405
timestamp 1666464484
transform 1 0 23352 0 -1 16464
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_413
timestamp 1666464484
transform 1 0 23800 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_417
timestamp 1666464484
transform 1 0 24024 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_419
timestamp 1666464484
transform 1 0 24136 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1666464484
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1666464484
transform 1 0 2576 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1666464484
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1666464484
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1666464484
transform 1 0 6552 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1666464484
transform 1 0 6720 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1666464484
transform 1 0 10304 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1666464484
transform 1 0 10528 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1666464484
transform 1 0 10696 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1666464484
transform 1 0 14280 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1666464484
transform 1 0 14504 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1666464484
transform 1 0 14672 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1666464484
transform 1 0 18256 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1666464484
transform 1 0 18480 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1666464484
transform 1 0 18648 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1666464484
transform 1 0 22232 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1666464484
transform 1 0 22456 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_392
timestamp 1666464484
transform 1 0 22624 0 1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_408
timestamp 1666464484
transform 1 0 23520 0 1 16464
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_416
timestamp 1666464484
transform 1 0 23968 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1666464484
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1666464484
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1666464484
transform 1 0 4592 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1666464484
transform 1 0 4760 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1666464484
transform 1 0 8344 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1666464484
transform 1 0 8568 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1666464484
transform 1 0 8736 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1666464484
transform 1 0 12320 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1666464484
transform 1 0 12544 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1666464484
transform 1 0 12712 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1666464484
transform 1 0 16296 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1666464484
transform 1 0 16520 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1666464484
transform 1 0 16688 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1666464484
transform 1 0 20272 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1666464484
transform 1 0 20496 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_357
timestamp 1666464484
transform 1 0 20664 0 -1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_389
timestamp 1666464484
transform 1 0 22456 0 -1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_405
timestamp 1666464484
transform 1 0 23352 0 -1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_413
timestamp 1666464484
transform 1 0 23800 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_417
timestamp 1666464484
transform 1 0 24024 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_419
timestamp 1666464484
transform 1 0 24136 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1666464484
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1666464484
transform 1 0 2576 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1666464484
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1666464484
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1666464484
transform 1 0 6552 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1666464484
transform 1 0 6720 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1666464484
transform 1 0 10304 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1666464484
transform 1 0 10528 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1666464484
transform 1 0 10696 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1666464484
transform 1 0 14280 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1666464484
transform 1 0 14504 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1666464484
transform 1 0 14672 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1666464484
transform 1 0 18256 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1666464484
transform 1 0 18480 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1666464484
transform 1 0 18648 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1666464484
transform 1 0 22232 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1666464484
transform 1 0 22456 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_392
timestamp 1666464484
transform 1 0 22624 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_408
timestamp 1666464484
transform 1 0 23520 0 1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_416
timestamp 1666464484
transform 1 0 23968 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1666464484
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_66
timestamp 1666464484
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1666464484
transform 1 0 4592 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1666464484
transform 1 0 4760 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1666464484
transform 1 0 8344 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1666464484
transform 1 0 8568 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1666464484
transform 1 0 8736 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1666464484
transform 1 0 12320 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1666464484
transform 1 0 12544 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1666464484
transform 1 0 12712 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1666464484
transform 1 0 16296 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1666464484
transform 1 0 16520 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1666464484
transform 1 0 16688 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1666464484
transform 1 0 20272 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1666464484
transform 1 0 20496 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_357
timestamp 1666464484
transform 1 0 20664 0 -1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_389
timestamp 1666464484
transform 1 0 22456 0 -1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_405
timestamp 1666464484
transform 1 0 23352 0 -1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_413
timestamp 1666464484
transform 1 0 23800 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_417
timestamp 1666464484
transform 1 0 24024 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_419
timestamp 1666464484
transform 1 0 24136 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1666464484
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1666464484
transform 1 0 2576 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1666464484
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1666464484
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1666464484
transform 1 0 6552 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_108
timestamp 1666464484
transform 1 0 6720 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_172
timestamp 1666464484
transform 1 0 10304 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1666464484
transform 1 0 10528 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_179
timestamp 1666464484
transform 1 0 10696 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_243
timestamp 1666464484
transform 1 0 14280 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1666464484
transform 1 0 14504 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_250
timestamp 1666464484
transform 1 0 14672 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_314
timestamp 1666464484
transform 1 0 18256 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1666464484
transform 1 0 18480 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_321
timestamp 1666464484
transform 1 0 18648 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_385
timestamp 1666464484
transform 1 0 22232 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_389
timestamp 1666464484
transform 1 0 22456 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_392
timestamp 1666464484
transform 1 0 22624 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_408
timestamp 1666464484
transform 1 0 23520 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_416
timestamp 1666464484
transform 1 0 23968 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_2
timestamp 1666464484
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_66
timestamp 1666464484
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_70
timestamp 1666464484
transform 1 0 4592 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_73
timestamp 1666464484
transform 1 0 4760 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_137
timestamp 1666464484
transform 1 0 8344 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1666464484
transform 1 0 8568 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_144
timestamp 1666464484
transform 1 0 8736 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_208
timestamp 1666464484
transform 1 0 12320 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1666464484
transform 1 0 12544 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1666464484
transform 1 0 12712 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_279
timestamp 1666464484
transform 1 0 16296 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1666464484
transform 1 0 16520 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_286
timestamp 1666464484
transform 1 0 16688 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_350
timestamp 1666464484
transform 1 0 20272 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1666464484
transform 1 0 20496 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_357
timestamp 1666464484
transform 1 0 20664 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_389
timestamp 1666464484
transform 1 0 22456 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_405
timestamp 1666464484
transform 1 0 23352 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_413
timestamp 1666464484
transform 1 0 23800 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_417
timestamp 1666464484
transform 1 0 24024 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_419
timestamp 1666464484
transform 1 0 24136 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_2
timestamp 1666464484
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1666464484
transform 1 0 2576 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_37
timestamp 1666464484
transform 1 0 2744 0 1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_101
timestamp 1666464484
transform 1 0 6328 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1666464484
transform 1 0 6552 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_108
timestamp 1666464484
transform 1 0 6720 0 1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_172
timestamp 1666464484
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1666464484
transform 1 0 10528 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_179
timestamp 1666464484
transform 1 0 10696 0 1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_243
timestamp 1666464484
transform 1 0 14280 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1666464484
transform 1 0 14504 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1666464484
transform 1 0 14672 0 1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_314
timestamp 1666464484
transform 1 0 18256 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1666464484
transform 1 0 18480 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_321
timestamp 1666464484
transform 1 0 18648 0 1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_385
timestamp 1666464484
transform 1 0 22232 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1666464484
transform 1 0 22456 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_392
timestamp 1666464484
transform 1 0 22624 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_408
timestamp 1666464484
transform 1 0 23520 0 1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_416
timestamp 1666464484
transform 1 0 23968 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_2
timestamp 1666464484
transform 1 0 784 0 -1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_66
timestamp 1666464484
transform 1 0 4368 0 -1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1666464484
transform 1 0 4592 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_73
timestamp 1666464484
transform 1 0 4760 0 -1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_137
timestamp 1666464484
transform 1 0 8344 0 -1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1666464484
transform 1 0 8568 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_144
timestamp 1666464484
transform 1 0 8736 0 -1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_208
timestamp 1666464484
transform 1 0 12320 0 -1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1666464484
transform 1 0 12544 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1666464484
transform 1 0 12712 0 -1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1666464484
transform 1 0 16296 0 -1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1666464484
transform 1 0 16520 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_286
timestamp 1666464484
transform 1 0 16688 0 -1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_350
timestamp 1666464484
transform 1 0 20272 0 -1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1666464484
transform 1 0 20496 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_357
timestamp 1666464484
transform 1 0 20664 0 -1 19600
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_389
timestamp 1666464484
transform 1 0 22456 0 -1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_405
timestamp 1666464484
transform 1 0 23352 0 -1 19600
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_413
timestamp 1666464484
transform 1 0 23800 0 -1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_417
timestamp 1666464484
transform 1 0 24024 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_419
timestamp 1666464484
transform 1 0 24136 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_2
timestamp 1666464484
transform 1 0 784 0 1 19600
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1666464484
transform 1 0 2576 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1666464484
transform 1 0 2744 0 1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1666464484
transform 1 0 6328 0 1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1666464484
transform 1 0 6552 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_108
timestamp 1666464484
transform 1 0 6720 0 1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_172
timestamp 1666464484
transform 1 0 10304 0 1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1666464484
transform 1 0 10528 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_179
timestamp 1666464484
transform 1 0 10696 0 1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_243
timestamp 1666464484
transform 1 0 14280 0 1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1666464484
transform 1 0 14504 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1666464484
transform 1 0 14672 0 1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_314
timestamp 1666464484
transform 1 0 18256 0 1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1666464484
transform 1 0 18480 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_321
timestamp 1666464484
transform 1 0 18648 0 1 19600
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_385
timestamp 1666464484
transform 1 0 22232 0 1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1666464484
transform 1 0 22456 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_392
timestamp 1666464484
transform 1 0 22624 0 1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_408
timestamp 1666464484
transform 1 0 23520 0 1 19600
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_416
timestamp 1666464484
transform 1 0 23968 0 1 19600
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_2
timestamp 1666464484
transform 1 0 784 0 -1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_66
timestamp 1666464484
transform 1 0 4368 0 -1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1666464484
transform 1 0 4592 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_73
timestamp 1666464484
transform 1 0 4760 0 -1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_137
timestamp 1666464484
transform 1 0 8344 0 -1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1666464484
transform 1 0 8568 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_144
timestamp 1666464484
transform 1 0 8736 0 -1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_208
timestamp 1666464484
transform 1 0 12320 0 -1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1666464484
transform 1 0 12544 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_215
timestamp 1666464484
transform 1 0 12712 0 -1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_279
timestamp 1666464484
transform 1 0 16296 0 -1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_283
timestamp 1666464484
transform 1 0 16520 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_286
timestamp 1666464484
transform 1 0 16688 0 -1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_350
timestamp 1666464484
transform 1 0 20272 0 -1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_354
timestamp 1666464484
transform 1 0 20496 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_357
timestamp 1666464484
transform 1 0 20664 0 -1 20384
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_389
timestamp 1666464484
transform 1 0 22456 0 -1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_405
timestamp 1666464484
transform 1 0 23352 0 -1 20384
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_413
timestamp 1666464484
transform 1 0 23800 0 -1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_417
timestamp 1666464484
transform 1 0 24024 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_419
timestamp 1666464484
transform 1 0 24136 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_2
timestamp 1666464484
transform 1 0 784 0 1 20384
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_34
timestamp 1666464484
transform 1 0 2576 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_37
timestamp 1666464484
transform 1 0 2744 0 1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_101
timestamp 1666464484
transform 1 0 6328 0 1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1666464484
transform 1 0 6552 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_108
timestamp 1666464484
transform 1 0 6720 0 1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_172
timestamp 1666464484
transform 1 0 10304 0 1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1666464484
transform 1 0 10528 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_179
timestamp 1666464484
transform 1 0 10696 0 1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_243
timestamp 1666464484
transform 1 0 14280 0 1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1666464484
transform 1 0 14504 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_250
timestamp 1666464484
transform 1 0 14672 0 1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_314
timestamp 1666464484
transform 1 0 18256 0 1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1666464484
transform 1 0 18480 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_321
timestamp 1666464484
transform 1 0 18648 0 1 20384
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_385
timestamp 1666464484
transform 1 0 22232 0 1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_389
timestamp 1666464484
transform 1 0 22456 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_392
timestamp 1666464484
transform 1 0 22624 0 1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_408
timestamp 1666464484
transform 1 0 23520 0 1 20384
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_416
timestamp 1666464484
transform 1 0 23968 0 1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_2
timestamp 1666464484
transform 1 0 784 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_7
timestamp 1666464484
transform 1 0 1064 0 -1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_73
timestamp 1666464484
transform 1 0 4760 0 -1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_137
timestamp 1666464484
transform 1 0 8344 0 -1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1666464484
transform 1 0 8568 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_144
timestamp 1666464484
transform 1 0 8736 0 -1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_208
timestamp 1666464484
transform 1 0 12320 0 -1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1666464484
transform 1 0 12544 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_215
timestamp 1666464484
transform 1 0 12712 0 -1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_279
timestamp 1666464484
transform 1 0 16296 0 -1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1666464484
transform 1 0 16520 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_286
timestamp 1666464484
transform 1 0 16688 0 -1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_350
timestamp 1666464484
transform 1 0 20272 0 -1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1666464484
transform 1 0 20496 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_357
timestamp 1666464484
transform 1 0 20664 0 -1 21168
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_389
timestamp 1666464484
transform 1 0 22456 0 -1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_405
timestamp 1666464484
transform 1 0 23352 0 -1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_413
timestamp 1666464484
transform 1 0 23800 0 -1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_417
timestamp 1666464484
transform 1 0 24024 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_419
timestamp 1666464484
transform 1 0 24136 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_2
timestamp 1666464484
transform 1 0 784 0 1 21168
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1666464484
transform 1 0 2576 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_37
timestamp 1666464484
transform 1 0 2744 0 1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_101
timestamp 1666464484
transform 1 0 6328 0 1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1666464484
transform 1 0 6552 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_108
timestamp 1666464484
transform 1 0 6720 0 1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_172
timestamp 1666464484
transform 1 0 10304 0 1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1666464484
transform 1 0 10528 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_179
timestamp 1666464484
transform 1 0 10696 0 1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_243
timestamp 1666464484
transform 1 0 14280 0 1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1666464484
transform 1 0 14504 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_250
timestamp 1666464484
transform 1 0 14672 0 1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_314
timestamp 1666464484
transform 1 0 18256 0 1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1666464484
transform 1 0 18480 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_321
timestamp 1666464484
transform 1 0 18648 0 1 21168
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_385
timestamp 1666464484
transform 1 0 22232 0 1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1666464484
transform 1 0 22456 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_392
timestamp 1666464484
transform 1 0 22624 0 1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_408
timestamp 1666464484
transform 1 0 23520 0 1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_416
timestamp 1666464484
transform 1 0 23968 0 1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_2
timestamp 1666464484
transform 1 0 784 0 -1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_66
timestamp 1666464484
transform 1 0 4368 0 -1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1666464484
transform 1 0 4592 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_73
timestamp 1666464484
transform 1 0 4760 0 -1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_137
timestamp 1666464484
transform 1 0 8344 0 -1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1666464484
transform 1 0 8568 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_144
timestamp 1666464484
transform 1 0 8736 0 -1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_208
timestamp 1666464484
transform 1 0 12320 0 -1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1666464484
transform 1 0 12544 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_215
timestamp 1666464484
transform 1 0 12712 0 -1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_279
timestamp 1666464484
transform 1 0 16296 0 -1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_283
timestamp 1666464484
transform 1 0 16520 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_286
timestamp 1666464484
transform 1 0 16688 0 -1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_350
timestamp 1666464484
transform 1 0 20272 0 -1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1666464484
transform 1 0 20496 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_357
timestamp 1666464484
transform 1 0 20664 0 -1 21952
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_389
timestamp 1666464484
transform 1 0 22456 0 -1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_405
timestamp 1666464484
transform 1 0 23352 0 -1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_413
timestamp 1666464484
transform 1 0 23800 0 -1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_417
timestamp 1666464484
transform 1 0 24024 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_419
timestamp 1666464484
transform 1 0 24136 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_2
timestamp 1666464484
transform 1 0 784 0 1 21952
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1666464484
transform 1 0 2576 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1666464484
transform 1 0 2744 0 1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1666464484
transform 1 0 6328 0 1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1666464484
transform 1 0 6552 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_108
timestamp 1666464484
transform 1 0 6720 0 1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_172
timestamp 1666464484
transform 1 0 10304 0 1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1666464484
transform 1 0 10528 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_179
timestamp 1666464484
transform 1 0 10696 0 1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_243
timestamp 1666464484
transform 1 0 14280 0 1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1666464484
transform 1 0 14504 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_250
timestamp 1666464484
transform 1 0 14672 0 1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_314
timestamp 1666464484
transform 1 0 18256 0 1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1666464484
transform 1 0 18480 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_321
timestamp 1666464484
transform 1 0 18648 0 1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_385
timestamp 1666464484
transform 1 0 22232 0 1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1666464484
transform 1 0 22456 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_392
timestamp 1666464484
transform 1 0 22624 0 1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_408
timestamp 1666464484
transform 1 0 23520 0 1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_416
timestamp 1666464484
transform 1 0 23968 0 1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_2
timestamp 1666464484
transform 1 0 784 0 -1 22736
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_66
timestamp 1666464484
transform 1 0 4368 0 -1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_70
timestamp 1666464484
transform 1 0 4592 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_73
timestamp 1666464484
transform 1 0 4760 0 -1 22736
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_137
timestamp 1666464484
transform 1 0 8344 0 -1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1666464484
transform 1 0 8568 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_144
timestamp 1666464484
transform 1 0 8736 0 -1 22736
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_208
timestamp 1666464484
transform 1 0 12320 0 -1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1666464484
transform 1 0 12544 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_215
timestamp 1666464484
transform 1 0 12712 0 -1 22736
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_279
timestamp 1666464484
transform 1 0 16296 0 -1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1666464484
transform 1 0 16520 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_286
timestamp 1666464484
transform 1 0 16688 0 -1 22736
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_350
timestamp 1666464484
transform 1 0 20272 0 -1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1666464484
transform 1 0 20496 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_357
timestamp 1666464484
transform 1 0 20664 0 -1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_389
timestamp 1666464484
transform 1 0 22456 0 -1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_405
timestamp 1666464484
transform 1 0 23352 0 -1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_413
timestamp 1666464484
transform 1 0 23800 0 -1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_417
timestamp 1666464484
transform 1 0 24024 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_419
timestamp 1666464484
transform 1 0 24136 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_2
timestamp 1666464484
transform 1 0 784 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1666464484
transform 1 0 2576 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_37
timestamp 1666464484
transform 1 0 2744 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_69
timestamp 1666464484
transform 1 0 4536 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_72
timestamp 1666464484
transform 1 0 4704 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_104
timestamp 1666464484
transform 1 0 6496 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_107
timestamp 1666464484
transform 1 0 6664 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_139
timestamp 1666464484
transform 1 0 8456 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_142
timestamp 1666464484
transform 1 0 8624 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_174
timestamp 1666464484
transform 1 0 10416 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_177
timestamp 1666464484
transform 1 0 10584 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_209
timestamp 1666464484
transform 1 0 12376 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_212
timestamp 1666464484
transform 1 0 12544 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_244
timestamp 1666464484
transform 1 0 14336 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_247
timestamp 1666464484
transform 1 0 14504 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_279
timestamp 1666464484
transform 1 0 16296 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_282
timestamp 1666464484
transform 1 0 16464 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_314
timestamp 1666464484
transform 1 0 18256 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_317
timestamp 1666464484
transform 1 0 18424 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_349
timestamp 1666464484
transform 1 0 20216 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_352
timestamp 1666464484
transform 1 0 20384 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_384
timestamp 1666464484
transform 1 0 22176 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_387
timestamp 1666464484
transform 1 0 22344 0 1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_419
timestamp 1666464484
transform 1 0 24136 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1666464484
transform -1 0 24304 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1666464484
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1666464484
transform -1 0 24304 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1666464484
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1666464484
transform -1 0 24304 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1666464484
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1666464484
transform -1 0 24304 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1666464484
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1666464484
transform -1 0 24304 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1666464484
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1666464484
transform -1 0 24304 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1666464484
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1666464484
transform -1 0 24304 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1666464484
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1666464484
transform -1 0 24304 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1666464484
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1666464484
transform -1 0 24304 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1666464484
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1666464484
transform -1 0 24304 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1666464484
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1666464484
transform -1 0 24304 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1666464484
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1666464484
transform -1 0 24304 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1666464484
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1666464484
transform -1 0 24304 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1666464484
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1666464484
transform -1 0 24304 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1666464484
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1666464484
transform -1 0 24304 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1666464484
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1666464484
transform -1 0 24304 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1666464484
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1666464484
transform -1 0 24304 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1666464484
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1666464484
transform -1 0 24304 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1666464484
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1666464484
transform -1 0 24304 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1666464484
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1666464484
transform -1 0 24304 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1666464484
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1666464484
transform -1 0 24304 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1666464484
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1666464484
transform -1 0 24304 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1666464484
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1666464484
transform -1 0 24304 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1666464484
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1666464484
transform -1 0 24304 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1666464484
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1666464484
transform -1 0 24304 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1666464484
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1666464484
transform -1 0 24304 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1666464484
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1666464484
transform -1 0 24304 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1666464484
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1666464484
transform -1 0 24304 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1666464484
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1666464484
transform -1 0 24304 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1666464484
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1666464484
transform -1 0 24304 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1666464484
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1666464484
transform -1 0 24304 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1666464484
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1666464484
transform -1 0 24304 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1666464484
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1666464484
transform -1 0 24304 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1666464484
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1666464484
transform -1 0 24304 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1666464484
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1666464484
transform -1 0 24304 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1666464484
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1666464484
transform -1 0 24304 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1666464484
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1666464484
transform -1 0 24304 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1666464484
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1666464484
transform -1 0 24304 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1666464484
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1666464484
transform -1 0 24304 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1666464484
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1666464484
transform -1 0 24304 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1666464484
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1666464484
transform -1 0 24304 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1666464484
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1666464484
transform -1 0 24304 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1666464484
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1666464484
transform -1 0 24304 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1666464484
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1666464484
transform -1 0 24304 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1666464484
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1666464484
transform -1 0 24304 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1666464484
transform 1 0 672 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1666464484
transform -1 0 24304 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1666464484
transform 1 0 672 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1666464484
transform -1 0 24304 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1666464484
transform 1 0 672 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1666464484
transform -1 0 24304 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1666464484
transform 1 0 672 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1666464484
transform -1 0 24304 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1666464484
transform 1 0 672 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1666464484
transform -1 0 24304 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1666464484
transform 1 0 672 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1666464484
transform -1 0 24304 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1666464484
transform 1 0 672 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1666464484
transform -1 0 24304 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1666464484
transform 1 0 672 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1666464484
transform -1 0 24304 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1666464484
transform 1 0 672 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1666464484
transform -1 0 24304 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1666464484
transform 1 0 672 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1666464484
transform -1 0 24304 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 2632 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1666464484
transform 1 0 4592 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1666464484
transform 1 0 6552 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1666464484
transform 1 0 8512 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1666464484
transform 1 0 10472 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1666464484
transform 1 0 12432 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1666464484
transform 1 0 14392 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1666464484
transform 1 0 16352 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1666464484
transform 1 0 18312 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1666464484
transform 1 0 20272 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1666464484
transform 1 0 22232 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1666464484
transform 1 0 4648 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1666464484
transform 1 0 8624 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1666464484
transform 1 0 12600 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1666464484
transform 1 0 16576 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1666464484
transform 1 0 20552 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1666464484
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1666464484
transform 1 0 6608 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1666464484
transform 1 0 10584 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1666464484
transform 1 0 14560 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1666464484
transform 1 0 18536 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1666464484
transform 1 0 22512 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1666464484
transform 1 0 4648 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1666464484
transform 1 0 8624 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1666464484
transform 1 0 12600 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1666464484
transform 1 0 16576 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1666464484
transform 1 0 20552 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1666464484
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1666464484
transform 1 0 6608 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1666464484
transform 1 0 10584 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1666464484
transform 1 0 14560 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1666464484
transform 1 0 18536 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1666464484
transform 1 0 22512 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1666464484
transform 1 0 4648 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1666464484
transform 1 0 8624 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1666464484
transform 1 0 12600 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1666464484
transform 1 0 16576 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1666464484
transform 1 0 20552 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1666464484
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1666464484
transform 1 0 6608 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1666464484
transform 1 0 10584 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1666464484
transform 1 0 14560 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1666464484
transform 1 0 18536 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1666464484
transform 1 0 22512 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1666464484
transform 1 0 4648 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1666464484
transform 1 0 8624 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1666464484
transform 1 0 12600 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1666464484
transform 1 0 16576 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1666464484
transform 1 0 20552 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1666464484
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1666464484
transform 1 0 6608 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1666464484
transform 1 0 10584 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1666464484
transform 1 0 14560 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1666464484
transform 1 0 18536 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1666464484
transform 1 0 22512 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1666464484
transform 1 0 4648 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1666464484
transform 1 0 8624 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1666464484
transform 1 0 12600 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1666464484
transform 1 0 16576 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1666464484
transform 1 0 20552 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1666464484
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1666464484
transform 1 0 6608 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1666464484
transform 1 0 10584 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1666464484
transform 1 0 14560 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1666464484
transform 1 0 18536 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1666464484
transform 1 0 22512 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1666464484
transform 1 0 4648 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1666464484
transform 1 0 8624 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1666464484
transform 1 0 12600 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1666464484
transform 1 0 16576 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1666464484
transform 1 0 20552 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1666464484
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1666464484
transform 1 0 6608 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1666464484
transform 1 0 10584 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1666464484
transform 1 0 14560 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1666464484
transform 1 0 18536 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1666464484
transform 1 0 22512 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1666464484
transform 1 0 4648 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1666464484
transform 1 0 8624 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1666464484
transform 1 0 12600 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1666464484
transform 1 0 16576 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1666464484
transform 1 0 20552 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1666464484
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1666464484
transform 1 0 6608 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1666464484
transform 1 0 10584 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1666464484
transform 1 0 14560 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1666464484
transform 1 0 18536 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1666464484
transform 1 0 22512 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1666464484
transform 1 0 4648 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1666464484
transform 1 0 8624 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1666464484
transform 1 0 12600 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1666464484
transform 1 0 16576 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1666464484
transform 1 0 20552 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1666464484
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1666464484
transform 1 0 6608 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1666464484
transform 1 0 10584 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1666464484
transform 1 0 14560 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1666464484
transform 1 0 18536 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1666464484
transform 1 0 22512 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1666464484
transform 1 0 4648 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1666464484
transform 1 0 8624 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1666464484
transform 1 0 12600 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1666464484
transform 1 0 16576 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1666464484
transform 1 0 20552 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1666464484
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1666464484
transform 1 0 6608 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1666464484
transform 1 0 10584 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1666464484
transform 1 0 14560 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1666464484
transform 1 0 18536 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1666464484
transform 1 0 22512 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1666464484
transform 1 0 4648 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1666464484
transform 1 0 8624 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1666464484
transform 1 0 12600 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1666464484
transform 1 0 16576 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1666464484
transform 1 0 20552 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1666464484
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1666464484
transform 1 0 6608 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1666464484
transform 1 0 10584 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1666464484
transform 1 0 14560 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1666464484
transform 1 0 18536 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1666464484
transform 1 0 22512 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1666464484
transform 1 0 4648 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1666464484
transform 1 0 8624 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1666464484
transform 1 0 12600 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1666464484
transform 1 0 16576 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1666464484
transform 1 0 20552 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1666464484
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1666464484
transform 1 0 6608 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1666464484
transform 1 0 10584 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1666464484
transform 1 0 14560 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1666464484
transform 1 0 18536 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1666464484
transform 1 0 22512 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1666464484
transform 1 0 4648 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1666464484
transform 1 0 8624 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1666464484
transform 1 0 12600 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1666464484
transform 1 0 16576 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1666464484
transform 1 0 20552 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1666464484
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1666464484
transform 1 0 6608 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1666464484
transform 1 0 10584 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1666464484
transform 1 0 14560 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1666464484
transform 1 0 18536 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1666464484
transform 1 0 22512 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1666464484
transform 1 0 4648 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1666464484
transform 1 0 8624 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1666464484
transform 1 0 12600 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1666464484
transform 1 0 16576 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1666464484
transform 1 0 20552 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1666464484
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1666464484
transform 1 0 6608 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1666464484
transform 1 0 10584 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1666464484
transform 1 0 14560 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1666464484
transform 1 0 18536 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1666464484
transform 1 0 22512 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1666464484
transform 1 0 4648 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1666464484
transform 1 0 8624 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1666464484
transform 1 0 12600 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1666464484
transform 1 0 16576 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1666464484
transform 1 0 20552 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1666464484
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1666464484
transform 1 0 6608 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1666464484
transform 1 0 10584 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1666464484
transform 1 0 14560 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1666464484
transform 1 0 18536 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1666464484
transform 1 0 22512 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1666464484
transform 1 0 4648 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1666464484
transform 1 0 8624 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1666464484
transform 1 0 12600 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1666464484
transform 1 0 16576 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1666464484
transform 1 0 20552 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1666464484
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1666464484
transform 1 0 6608 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1666464484
transform 1 0 10584 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1666464484
transform 1 0 14560 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1666464484
transform 1 0 18536 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1666464484
transform 1 0 22512 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1666464484
transform 1 0 4648 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1666464484
transform 1 0 8624 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1666464484
transform 1 0 12600 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1666464484
transform 1 0 16576 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1666464484
transform 1 0 20552 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1666464484
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1666464484
transform 1 0 6608 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1666464484
transform 1 0 10584 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1666464484
transform 1 0 14560 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1666464484
transform 1 0 18536 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1666464484
transform 1 0 22512 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1666464484
transform 1 0 4648 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1666464484
transform 1 0 8624 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1666464484
transform 1 0 12600 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1666464484
transform 1 0 16576 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1666464484
transform 1 0 20552 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1666464484
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1666464484
transform 1 0 6608 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1666464484
transform 1 0 10584 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1666464484
transform 1 0 14560 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1666464484
transform 1 0 18536 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1666464484
transform 1 0 22512 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1666464484
transform 1 0 4648 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1666464484
transform 1 0 8624 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1666464484
transform 1 0 12600 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1666464484
transform 1 0 16576 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1666464484
transform 1 0 20552 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1666464484
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1666464484
transform 1 0 6608 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1666464484
transform 1 0 10584 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1666464484
transform 1 0 14560 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1666464484
transform 1 0 18536 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1666464484
transform 1 0 22512 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1666464484
transform 1 0 4648 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1666464484
transform 1 0 8624 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1666464484
transform 1 0 12600 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1666464484
transform 1 0 16576 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1666464484
transform 1 0 20552 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1666464484
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1666464484
transform 1 0 6608 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1666464484
transform 1 0 10584 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1666464484
transform 1 0 14560 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1666464484
transform 1 0 18536 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1666464484
transform 1 0 22512 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1666464484
transform 1 0 4648 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1666464484
transform 1 0 8624 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1666464484
transform 1 0 12600 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1666464484
transform 1 0 16576 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1666464484
transform 1 0 20552 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1666464484
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1666464484
transform 1 0 6608 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1666464484
transform 1 0 10584 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1666464484
transform 1 0 14560 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1666464484
transform 1 0 18536 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1666464484
transform 1 0 22512 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1666464484
transform 1 0 4648 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1666464484
transform 1 0 8624 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1666464484
transform 1 0 12600 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1666464484
transform 1 0 16576 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1666464484
transform 1 0 20552 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1666464484
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1666464484
transform 1 0 6608 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1666464484
transform 1 0 10584 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1666464484
transform 1 0 14560 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1666464484
transform 1 0 18536 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1666464484
transform 1 0 22512 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1666464484
transform 1 0 4648 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1666464484
transform 1 0 8624 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1666464484
transform 1 0 12600 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1666464484
transform 1 0 16576 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1666464484
transform 1 0 20552 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1666464484
transform 1 0 2632 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1666464484
transform 1 0 6608 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1666464484
transform 1 0 10584 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1666464484
transform 1 0 14560 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1666464484
transform 1 0 18536 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1666464484
transform 1 0 22512 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1666464484
transform 1 0 4648 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1666464484
transform 1 0 8624 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1666464484
transform 1 0 12600 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1666464484
transform 1 0 16576 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1666464484
transform 1 0 20552 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1666464484
transform 1 0 2632 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1666464484
transform 1 0 6608 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1666464484
transform 1 0 10584 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1666464484
transform 1 0 14560 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1666464484
transform 1 0 18536 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1666464484
transform 1 0 22512 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1666464484
transform 1 0 4648 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1666464484
transform 1 0 8624 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1666464484
transform 1 0 12600 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1666464484
transform 1 0 16576 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1666464484
transform 1 0 20552 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1666464484
transform 1 0 2632 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1666464484
transform 1 0 6608 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1666464484
transform 1 0 10584 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1666464484
transform 1 0 14560 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1666464484
transform 1 0 18536 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1666464484
transform 1 0 22512 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1666464484
transform 1 0 4648 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1666464484
transform 1 0 8624 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1666464484
transform 1 0 12600 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1666464484
transform 1 0 16576 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1666464484
transform 1 0 20552 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1666464484
transform 1 0 2632 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1666464484
transform 1 0 6608 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1666464484
transform 1 0 10584 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1666464484
transform 1 0 14560 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1666464484
transform 1 0 18536 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1666464484
transform 1 0 22512 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1666464484
transform 1 0 4648 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1666464484
transform 1 0 8624 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1666464484
transform 1 0 12600 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1666464484
transform 1 0 16576 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1666464484
transform 1 0 20552 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1666464484
transform 1 0 2632 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1666464484
transform 1 0 6608 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1666464484
transform 1 0 10584 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1666464484
transform 1 0 14560 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1666464484
transform 1 0 18536 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1666464484
transform 1 0 22512 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1666464484
transform 1 0 4648 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1666464484
transform 1 0 8624 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1666464484
transform 1 0 12600 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1666464484
transform 1 0 16576 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1666464484
transform 1 0 20552 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1666464484
transform 1 0 2632 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1666464484
transform 1 0 4592 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1666464484
transform 1 0 6552 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1666464484
transform 1 0 8512 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1666464484
transform 1 0 10472 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1666464484
transform 1 0 12432 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1666464484
transform 1 0 14392 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1666464484
transform 1 0 16352 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1666464484
transform 1 0 18312 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1666464484
transform 1 0 20272 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1666464484
transform 1 0 22232 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 12208 0 1 5488
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 11984 0 -1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 11816 0 1 4704
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_core_clock dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform 1 0 12768 0 -1 5488
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_core_clock
timestamp 1666464484
transform -1 0 12320 0 -1 3920
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_core_clock
timestamp 1666464484
transform -1 0 16128 0 -1 6272
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  clock_source_sel_3 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 1064 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  clock_source_sel_4
timestamp 1666464484
transform -1 0 1064 0 -1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1666464484
transform -1 0 19096 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output2
timestamp 1666464484
transform -1 0 1176 0 -1 4704
box -43 -43 379 435
<< labels >>
flabel metal3 s -480 4116 240 4228 0 FreeSans 448 0 0 0 clock_out_a
port 0 nsew signal tristate
flabel metal3 s -480 12404 240 12516 0 FreeSans 448 0 0 0 clock_out_b
port 1 nsew signal tristate
flabel metal3 s -480 20692 240 20804 0 FreeSans 448 0 0 0 clock_out_c
port 2 nsew signal tristate
flabel metal2 s 6188 -480 6300 240 0 FreeSans 448 90 0 0 core_clock
port 3 nsew signal input
flabel metal3 s 24760 12404 25480 12516 0 FreeSans 448 0 0 0 io_clock
port 4 nsew signal input
flabel metal2 s 18676 -480 18788 240 0 FreeSans 448 90 0 0 la_oenb
port 5 nsew signal input
flabel metal4 s 1017 1538 1327 23158 0 FreeSans 1280 90 0 0 vccd1
port 6 nsew power bidirectional
flabel metal4 s 19017 1538 19327 23158 0 FreeSans 1280 90 0 0 vccd1
port 6 nsew power bidirectional
flabel metal4 s 2877 1538 3187 23158 0 FreeSans 1280 90 0 0 vssd1
port 7 nsew ground bidirectional
flabel metal4 s 20877 1538 21187 23158 0 FreeSans 1280 90 0 0 vssd1
port 7 nsew ground bidirectional
rlabel metal1 12488 23128 12488 23128 0 vccd1
rlabel metal1 12488 22736 12488 22736 0 vssd1
rlabel metal2 11900 5488 11900 5488 0 _0_
rlabel metal2 12348 3724 12348 3724 0 clknet_0_core_clock
rlabel metal3 11396 4900 11396 4900 0 clknet_1_0__leaf_core_clock
rlabel metal2 12908 5824 12908 5824 0 clknet_1_1__leaf_core_clock
rlabel metal3 567 4172 567 4172 0 clock_out_a
rlabel metal2 12852 5264 12852 5264 0 core_clock
rlabel metal3 23513 12460 23513 12460 0 io_clock
rlabel metal2 18648 1708 18648 1708 0 la_oenb
rlabel metal2 12292 4816 12292 4816 0 net1
rlabel metal3 1232 4508 1232 4508 0 net2
rlabel metal3 567 12516 567 12516 0 net3
rlabel metal3 567 20804 567 20804 0 net4
rlabel metal2 12852 5544 12852 5544 0 sel_reg
<< properties >>
string FIXED_BBOX 0 0 25000 25000
<< end >>
