// This is the unpowered netlist.
module controller_core (clock,
    io_control_trigger_in,
    io_control_trigger_oeb,
    io_latch_data_in,
    io_latch_data_oeb,
    io_reset_n_in,
    io_reset_n_oeb,
    io_update_cycle_complete_oeb,
    io_update_cycle_complete_out,
    output_active_left,
    output_active_right,
    spi_data_clock,
    clock_out,
    col_select_left,
    col_select_right,
    data_out_left,
    data_out_right,
    inverter_select,
    io_driver_io_oeb,
    la_data_in,
    la_oenb,
    mem_address_left,
    mem_address_right,
    mem_write_n,
    row_col_select,
    row_select_left,
    row_select_right,
    spi_data);
 input clock;
 input io_control_trigger_in;
 output io_control_trigger_oeb;
 input io_latch_data_in;
 output io_latch_data_oeb;
 input io_reset_n_in;
 output io_reset_n_oeb;
 output io_update_cycle_complete_oeb;
 output io_update_cycle_complete_out;
 output output_active_left;
 output output_active_right;
 input spi_data_clock;
 output [9:0] clock_out;
 output [5:0] col_select_left;
 output [5:0] col_select_right;
 output [15:0] data_out_left;
 output [15:0] data_out_right;
 output [9:0] inverter_select;
 output [19:0] io_driver_io_oeb;
 input [17:0] la_data_in;
 input [17:0] la_oenb;
 output [9:0] mem_address_left;
 output [9:0] mem_address_right;
 output [9:0] mem_write_n;
 output [9:0] row_col_select;
 output [5:0] row_select_left;
 output [5:0] row_select_right;
 input [31:0] spi_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire control_trigger;
 wire \control_trigger_sync[0] ;
 wire \control_trigger_sync[1] ;
 wire latch_data;
 wire \latch_data_sync[0] ;
 wire \latch_data_sync[1] ;
 wire reset_n;
 wire \reset_n_sync[0] ;
 wire \reset_n_sync[1] ;
 wire \spi_data_crossing[0].A ;
 wire \spi_data_crossing[0].data_sync ;
 wire \spi_data_crossing[10].A ;
 wire \spi_data_crossing[10].data_sync ;
 wire \spi_data_crossing[11].A ;
 wire \spi_data_crossing[11].data_sync ;
 wire \spi_data_crossing[12].A ;
 wire \spi_data_crossing[12].data_sync ;
 wire \spi_data_crossing[13].A ;
 wire \spi_data_crossing[13].data_sync ;
 wire \spi_data_crossing[14].A ;
 wire \spi_data_crossing[14].data_sync ;
 wire \spi_data_crossing[15].A ;
 wire \spi_data_crossing[15].data_sync ;
 wire \spi_data_crossing[16].A ;
 wire \spi_data_crossing[16].data_sync ;
 wire \spi_data_crossing[17].A ;
 wire \spi_data_crossing[17].data_sync ;
 wire \spi_data_crossing[18].A ;
 wire \spi_data_crossing[18].data_sync ;
 wire \spi_data_crossing[19].A ;
 wire \spi_data_crossing[19].data_sync ;
 wire \spi_data_crossing[1].A ;
 wire \spi_data_crossing[1].data_sync ;
 wire \spi_data_crossing[20].A ;
 wire \spi_data_crossing[20].data_sync ;
 wire \spi_data_crossing[21].A ;
 wire \spi_data_crossing[21].data_sync ;
 wire \spi_data_crossing[22].A ;
 wire \spi_data_crossing[22].data_sync ;
 wire \spi_data_crossing[23].A ;
 wire \spi_data_crossing[23].data_sync ;
 wire \spi_data_crossing[24].A ;
 wire \spi_data_crossing[24].data_sync ;
 wire \spi_data_crossing[25].A ;
 wire \spi_data_crossing[25].data_sync ;
 wire \spi_data_crossing[26].A ;
 wire \spi_data_crossing[26].data_sync ;
 wire \spi_data_crossing[27].A ;
 wire \spi_data_crossing[27].data_sync ;
 wire \spi_data_crossing[28].A ;
 wire \spi_data_crossing[28].data_sync ;
 wire \spi_data_crossing[29].A ;
 wire \spi_data_crossing[29].data_sync ;
 wire \spi_data_crossing[2].A ;
 wire \spi_data_crossing[2].data_sync ;
 wire \spi_data_crossing[30].A ;
 wire \spi_data_crossing[30].data_sync ;
 wire \spi_data_crossing[31].A ;
 wire \spi_data_crossing[31].data_sync ;
 wire \spi_data_crossing[3].A ;
 wire \spi_data_crossing[3].data_sync ;
 wire \spi_data_crossing[4].A ;
 wire \spi_data_crossing[4].data_sync ;
 wire \spi_data_crossing[5].A ;
 wire \spi_data_crossing[5].data_sync ;
 wire \spi_data_crossing[6].A ;
 wire \spi_data_crossing[6].data_sync ;
 wire \spi_data_crossing[7].A ;
 wire \spi_data_crossing[7].data_sync ;
 wire \spi_data_crossing[8].A ;
 wire \spi_data_crossing[8].data_sync ;
 wire \spi_data_crossing[9].A ;
 wire \spi_data_crossing[9].data_sync ;
 wire \u0.cmd[0] ;
 wire \u0.cmd[10] ;
 wire \u0.cmd[11] ;
 wire \u0.cmd[12] ;
 wire \u0.cmd[13] ;
 wire \u0.cmd[14] ;
 wire \u0.cmd[15] ;
 wire \u0.cmd[16] ;
 wire \u0.cmd[17] ;
 wire \u0.cmd[18] ;
 wire \u0.cmd[19] ;
 wire \u0.cmd[1] ;
 wire \u0.cmd[20] ;
 wire \u0.cmd[21] ;
 wire \u0.cmd[22] ;
 wire \u0.cmd[23] ;
 wire \u0.cmd[24] ;
 wire \u0.cmd[25] ;
 wire \u0.cmd[26] ;
 wire \u0.cmd[27] ;
 wire \u0.cmd[28] ;
 wire \u0.cmd[29] ;
 wire \u0.cmd[2] ;
 wire \u0.cmd[30] ;
 wire \u0.cmd[31] ;
 wire \u0.cmd[3] ;
 wire \u0.cmd[4] ;
 wire \u0.cmd[5] ;
 wire \u0.cmd[6] ;
 wire \u0.cmd[7] ;
 wire \u0.cmd[8] ;
 wire \u0.cmd[9] ;
 wire \u0.latch_cmd ;
 wire \u0.mem_write_n[0] ;
 wire \u0.mem_write_n[1] ;
 wire \u0.mem_write_n[2] ;
 wire \u0.mem_write_n[3] ;
 wire \u0.mem_write_n[4] ;
 wire \u0.mem_write_n[5] ;
 wire \u0.mem_write_n[6] ;
 wire \u0.mem_write_n[7] ;
 wire \u0.mem_write_n[8] ;
 wire \u0.mem_write_n[9] ;
 wire \u0.run_state[0] ;
 wire \u0.run_state[1] ;
 wire \u0.run_state[2] ;
 wire \u0.run_state[3] ;
 wire \u0.run_state[4] ;
 wire \u0.run_state[5] ;
 wire \u0.run_state[6] ;
 wire \u0.timer_enable ;
 wire \u0.u11.impulse_gen[0] ;
 wire \u0.u11.impulse_gen[1] ;
 wire \u0.update_cmd ;
 wire \u0.write_config_n ;
 wire \u1.ccr0[0] ;
 wire \u1.ccr0[10] ;
 wire \u1.ccr0[11] ;
 wire \u1.ccr0[12] ;
 wire \u1.ccr0[13] ;
 wire \u1.ccr0[14] ;
 wire \u1.ccr0[15] ;
 wire \u1.ccr0[16] ;
 wire \u1.ccr0[17] ;
 wire \u1.ccr0[18] ;
 wire \u1.ccr0[19] ;
 wire \u1.ccr0[1] ;
 wire \u1.ccr0[20] ;
 wire \u1.ccr0[21] ;
 wire \u1.ccr0[22] ;
 wire \u1.ccr0[23] ;
 wire \u1.ccr0[24] ;
 wire \u1.ccr0[25] ;
 wire \u1.ccr0[26] ;
 wire \u1.ccr0[27] ;
 wire \u1.ccr0[28] ;
 wire \u1.ccr0[29] ;
 wire \u1.ccr0[2] ;
 wire \u1.ccr0[30] ;
 wire \u1.ccr0[31] ;
 wire \u1.ccr0[3] ;
 wire \u1.ccr0[4] ;
 wire \u1.ccr0[5] ;
 wire \u1.ccr0[6] ;
 wire \u1.ccr0[7] ;
 wire \u1.ccr0[8] ;
 wire \u1.ccr0[9] ;
 wire \u1.ccr1[0] ;
 wire \u1.ccr1[10] ;
 wire \u1.ccr1[11] ;
 wire \u1.ccr1[12] ;
 wire \u1.ccr1[13] ;
 wire \u1.ccr1[14] ;
 wire \u1.ccr1[15] ;
 wire \u1.ccr1[16] ;
 wire \u1.ccr1[17] ;
 wire \u1.ccr1[18] ;
 wire \u1.ccr1[19] ;
 wire \u1.ccr1[1] ;
 wire \u1.ccr1[20] ;
 wire \u1.ccr1[21] ;
 wire \u1.ccr1[22] ;
 wire \u1.ccr1[23] ;
 wire \u1.ccr1[24] ;
 wire \u1.ccr1[25] ;
 wire \u1.ccr1[26] ;
 wire \u1.ccr1[27] ;
 wire \u1.ccr1[28] ;
 wire \u1.ccr1[29] ;
 wire \u1.ccr1[2] ;
 wire \u1.ccr1[30] ;
 wire \u1.ccr1[31] ;
 wire \u1.ccr1[3] ;
 wire \u1.ccr1[4] ;
 wire \u1.ccr1[5] ;
 wire \u1.ccr1[6] ;
 wire \u1.ccr1[7] ;
 wire \u1.ccr1[8] ;
 wire \u1.ccr1[9] ;
 wire \u1.ccr1_flag ;
 wire \u1.col_limit[0] ;
 wire \u1.col_limit[1] ;
 wire \u1.col_limit[2] ;
 wire \u1.col_limit[3] ;
 wire \u1.col_limit[4] ;
 wire \u1.col_limit[5] ;
 wire \u1.col_limit[6] ;
 wire \u1.col_sel[0] ;
 wire \u1.col_sel[1] ;
 wire \u1.col_sel[2] ;
 wire \u1.col_sel[3] ;
 wire \u1.col_sel[4] ;
 wire \u1.col_sel[5] ;
 wire \u1.col_sel[6] ;
 wire \u1.inverter_select[0] ;
 wire \u1.inverter_select[1] ;
 wire \u1.inverter_select[2] ;
 wire \u1.inverter_select[3] ;
 wire \u1.inverter_select[4] ;
 wire \u1.inverter_select[5] ;
 wire \u1.inverter_select[6] ;
 wire \u1.inverter_select[7] ;
 wire \u1.inverter_select[8] ;
 wire \u1.inverter_select[9] ;
 wire \u1.ordering_complete[0] ;
 wire \u1.ordering_complete[10] ;
 wire \u1.ordering_complete[11] ;
 wire \u1.ordering_complete[12] ;
 wire \u1.ordering_complete[13] ;
 wire \u1.ordering_complete[14] ;
 wire \u1.ordering_complete[15] ;
 wire \u1.ordering_complete[16] ;
 wire \u1.ordering_complete[17] ;
 wire \u1.ordering_complete[18] ;
 wire \u1.ordering_complete[19] ;
 wire \u1.ordering_complete[1] ;
 wire \u1.ordering_complete[20] ;
 wire \u1.ordering_complete[21] ;
 wire \u1.ordering_complete[22] ;
 wire \u1.ordering_complete[23] ;
 wire \u1.ordering_complete[24] ;
 wire \u1.ordering_complete[25] ;
 wire \u1.ordering_complete[26] ;
 wire \u1.ordering_complete[27] ;
 wire \u1.ordering_complete[28] ;
 wire \u1.ordering_complete[29] ;
 wire \u1.ordering_complete[2] ;
 wire \u1.ordering_complete[30] ;
 wire \u1.ordering_complete[31] ;
 wire \u1.ordering_complete[3] ;
 wire \u1.ordering_complete[4] ;
 wire \u1.ordering_complete[5] ;
 wire \u1.ordering_complete[6] ;
 wire \u1.ordering_complete[7] ;
 wire \u1.ordering_complete[8] ;
 wire \u1.ordering_complete[9] ;
 wire \u1.ordering_timer[0] ;
 wire \u1.ordering_timer[10] ;
 wire \u1.ordering_timer[11] ;
 wire \u1.ordering_timer[12] ;
 wire \u1.ordering_timer[13] ;
 wire \u1.ordering_timer[14] ;
 wire \u1.ordering_timer[15] ;
 wire \u1.ordering_timer[16] ;
 wire \u1.ordering_timer[17] ;
 wire \u1.ordering_timer[18] ;
 wire \u1.ordering_timer[19] ;
 wire \u1.ordering_timer[1] ;
 wire \u1.ordering_timer[20] ;
 wire \u1.ordering_timer[21] ;
 wire \u1.ordering_timer[22] ;
 wire \u1.ordering_timer[23] ;
 wire \u1.ordering_timer[24] ;
 wire \u1.ordering_timer[25] ;
 wire \u1.ordering_timer[26] ;
 wire \u1.ordering_timer[27] ;
 wire \u1.ordering_timer[28] ;
 wire \u1.ordering_timer[29] ;
 wire \u1.ordering_timer[2] ;
 wire \u1.ordering_timer[30] ;
 wire \u1.ordering_timer[31] ;
 wire \u1.ordering_timer[3] ;
 wire \u1.ordering_timer[4] ;
 wire \u1.ordering_timer[5] ;
 wire \u1.ordering_timer[6] ;
 wire \u1.ordering_timer[7] ;
 wire \u1.ordering_timer[8] ;
 wire \u1.ordering_timer[9] ;
 wire \u1.output_active ;
 wire \u1.row_col_select[0] ;
 wire \u1.row_col_select[1] ;
 wire \u1.row_col_select[2] ;
 wire \u1.row_col_select[3] ;
 wire \u1.row_col_select[4] ;
 wire \u1.row_col_select[5] ;
 wire \u1.row_col_select[6] ;
 wire \u1.row_col_select[7] ;
 wire \u1.row_col_select[8] ;
 wire \u1.row_col_select[9] ;
 wire \u1.row_limit[0] ;
 wire \u1.row_limit[1] ;
 wire \u1.row_limit[2] ;
 wire \u1.row_limit[3] ;
 wire \u1.row_limit[4] ;
 wire \u1.row_limit[5] ;
 wire \u1.row_limit[6] ;
 wire \u1.row_sel[0] ;
 wire \u1.row_sel[1] ;
 wire \u1.row_sel[2] ;
 wire \u1.row_sel[3] ;
 wire \u1.row_sel[4] ;
 wire \u1.row_sel[5] ;
 wire \u1.row_sel[6] ;
 wire \u1.timer[0] ;
 wire \u1.timer[10] ;
 wire \u1.timer[11] ;
 wire \u1.timer[12] ;
 wire \u1.timer[13] ;
 wire \u1.timer[14] ;
 wire \u1.timer[15] ;
 wire \u1.timer[16] ;
 wire \u1.timer[17] ;
 wire \u1.timer[18] ;
 wire \u1.timer[19] ;
 wire \u1.timer[1] ;
 wire \u1.timer[20] ;
 wire \u1.timer[21] ;
 wire \u1.timer[22] ;
 wire \u1.timer[23] ;
 wire \u1.timer[24] ;
 wire \u1.timer[25] ;
 wire \u1.timer[26] ;
 wire \u1.timer[27] ;
 wire \u1.timer[28] ;
 wire \u1.timer[29] ;
 wire \u1.timer[2] ;
 wire \u1.timer[30] ;
 wire \u1.timer[31] ;
 wire \u1.timer[3] ;
 wire \u1.timer[4] ;
 wire \u1.timer[5] ;
 wire \u1.timer[6] ;
 wire \u1.timer[7] ;
 wire \u1.timer[8] ;
 wire \u1.timer[9] ;
 wire \u1.u1.impulse_gen[0] ;
 wire \u1.u1.impulse_gen[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire clknet_leaf_0_clock;
 wire clknet_leaf_1_clock;
 wire clknet_leaf_2_clock;
 wire clknet_leaf_3_clock;
 wire clknet_leaf_4_clock;
 wire clknet_leaf_5_clock;
 wire clknet_leaf_6_clock;
 wire clknet_leaf_7_clock;
 wire clknet_leaf_8_clock;
 wire clknet_leaf_9_clock;
 wire clknet_leaf_10_clock;
 wire clknet_leaf_11_clock;
 wire clknet_leaf_12_clock;
 wire clknet_leaf_13_clock;
 wire clknet_leaf_14_clock;
 wire clknet_leaf_15_clock;
 wire clknet_leaf_16_clock;
 wire clknet_leaf_17_clock;
 wire clknet_leaf_18_clock;
 wire clknet_leaf_19_clock;
 wire clknet_leaf_20_clock;
 wire clknet_leaf_21_clock;
 wire clknet_leaf_22_clock;
 wire clknet_leaf_23_clock;
 wire clknet_leaf_24_clock;
 wire clknet_leaf_25_clock;
 wire clknet_leaf_26_clock;
 wire clknet_leaf_27_clock;
 wire clknet_leaf_28_clock;
 wire clknet_leaf_29_clock;
 wire clknet_leaf_30_clock;
 wire clknet_leaf_31_clock;
 wire clknet_leaf_32_clock;
 wire clknet_leaf_33_clock;
 wire clknet_leaf_34_clock;
 wire clknet_leaf_35_clock;
 wire clknet_leaf_36_clock;
 wire clknet_leaf_37_clock;
 wire clknet_leaf_38_clock;
 wire clknet_0_clock;
 wire clknet_2_0__leaf_clock;
 wire clknet_2_1__leaf_clock;
 wire clknet_2_2__leaf_clock;
 wire clknet_2_3__leaf_clock;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1415_ (.I(\u0.cmd[31] ),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1416_ (.A1(\reset_n_sync[1] ),
    .A2(\reset_n_sync[0] ),
    .A3(reset_n),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1417_ (.I(_1041_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1418_ (.A1(_1040_),
    .A2(\u0.cmd[30] ),
    .A3(_1042_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1419_ (.A1(\control_trigger_sync[0] ),
    .A2(control_trigger),
    .A3(\control_trigger_sync[1] ),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1420_ (.A1(\u0.cmd[26] ),
    .A2(_1044_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1421_ (.I(\u1.ordering_timer[23] ),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1422_ (.I(\u1.ordering_timer[22] ),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1423_ (.A1(_1046_),
    .A2(\u1.ordering_complete[23] ),
    .B1(_1047_),
    .B2(\u1.ordering_complete[22] ),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1424_ (.I(\u1.ordering_timer[21] ),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1425_ (.I(\u1.ordering_timer[20] ),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1426_ (.A1(_1049_),
    .A2(\u1.ordering_complete[21] ),
    .B1(_1050_),
    .B2(\u1.ordering_complete[20] ),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1427_ (.A1(_1048_),
    .A2(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1428_ (.A1(_1047_),
    .A2(\u1.ordering_complete[22] ),
    .B1(_1049_),
    .B2(\u1.ordering_complete[21] ),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1429_ (.I(\u1.ordering_complete[23] ),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1430_ (.A1(\u1.ordering_timer[23] ),
    .A2(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1431_ (.A1(_1050_),
    .A2(\u1.ordering_complete[20] ),
    .B(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1432_ (.A1(_1052_),
    .A2(_1053_),
    .A3(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1433_ (.I(\u1.ordering_complete[19] ),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1434_ (.I(\u1.ordering_timer[16] ),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1435_ (.I(\u1.ordering_complete[16] ),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1436_ (.I(\u1.ordering_complete[17] ),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1437_ (.A1(\u1.ordering_timer[17] ),
    .A2(_1061_),
    .B1(\u1.ordering_timer[16] ),
    .B2(_1060_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1438_ (.A1(\u1.ordering_timer[19] ),
    .A2(_1058_),
    .B1(_1059_),
    .B2(_1060_),
    .C(_1062_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1439_ (.I(\u1.ordering_timer[19] ),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1440_ (.I(\u1.ordering_timer[18] ),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1441_ (.A1(_1064_),
    .A2(\u1.ordering_complete[19] ),
    .B1(_1065_),
    .B2(\u1.ordering_complete[18] ),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1442_ (.I(\u1.ordering_complete[18] ),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1443_ (.I(\u1.ordering_timer[17] ),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1444_ (.A1(\u1.ordering_timer[18] ),
    .A2(_1067_),
    .B1(_1068_),
    .B2(_1061_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1445_ (.A1(_1057_),
    .A2(_1063_),
    .A3(_1066_),
    .A4(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1446_ (.I(\u1.ordering_timer[28] ),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1447_ (.I(\u1.ordering_timer[27] ),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1448_ (.I(\u1.ordering_complete[31] ),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1449_ (.A1(\u1.ordering_timer[31] ),
    .A2(_1073_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1450_ (.A1(_1071_),
    .A2(\u1.ordering_complete[28] ),
    .B1(_1072_),
    .B2(\u1.ordering_complete[27] ),
    .C(_1074_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1451_ (.I(\u1.ordering_timer[29] ),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1452_ (.A1(_1076_),
    .A2(\u1.ordering_complete[29] ),
    .B1(_1071_),
    .B2(\u1.ordering_complete[28] ),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1453_ (.I(\u1.ordering_complete[30] ),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1454_ (.I(\u1.ordering_complete[29] ),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1455_ (.A1(\u1.ordering_timer[30] ),
    .A2(_1078_),
    .B1(\u1.ordering_timer[29] ),
    .B2(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1456_ (.A1(_1077_),
    .A2(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1457_ (.I(\u1.ordering_timer[30] ),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1458_ (.A1(\u1.ordering_timer[31] ),
    .A2(_1073_),
    .B1(_1082_),
    .B2(_1078_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1459_ (.A1(_1075_),
    .A2(_1081_),
    .A3(_1083_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1460_ (.I(\u1.ordering_timer[24] ),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1461_ (.I(\u1.ordering_complete[24] ),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1462_ (.I(\u1.ordering_timer[26] ),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1463_ (.I(\u1.ordering_timer[25] ),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1464_ (.A1(_1087_),
    .A2(\u1.ordering_complete[26] ),
    .B1(_1088_),
    .B2(\u1.ordering_complete[25] ),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1465_ (.A1(_1085_),
    .A2(_1086_),
    .B(_1089_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1466_ (.A1(\u1.ordering_timer[24] ),
    .A2(_1086_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1467_ (.A1(_1088_),
    .A2(\u1.ordering_complete[25] ),
    .B(_1091_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1468_ (.I(_1072_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1469_ (.A1(_1093_),
    .A2(\u1.ordering_complete[27] ),
    .B1(_1087_),
    .B2(\u1.ordering_complete[26] ),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1470_ (.A1(_1084_),
    .A2(_1090_),
    .A3(_1092_),
    .A4(_1094_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1471_ (.I(\u1.ordering_timer[15] ),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1472_ (.I(\u1.ordering_complete[15] ),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1473_ (.I(\u1.ordering_complete[14] ),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1474_ (.A1(_1096_),
    .A2(_1097_),
    .B1(\u1.ordering_timer[14] ),
    .B2(_1098_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1475_ (.I(\u1.ordering_timer[14] ),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1476_ (.I(\u1.ordering_timer[13] ),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1477_ (.A1(_1100_),
    .A2(\u1.ordering_complete[14] ),
    .B1(_1101_),
    .B2(\u1.ordering_complete[13] ),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1478_ (.I(\u1.ordering_timer[12] ),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1479_ (.I(\u1.ordering_complete[11] ),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1480_ (.A1(\u1.ordering_timer[15] ),
    .A2(_1097_),
    .B1(\u1.ordering_timer[11] ),
    .B2(_1104_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1481_ (.A1(_1101_),
    .A2(\u1.ordering_complete[13] ),
    .B1(_1103_),
    .B2(\u1.ordering_complete[12] ),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1482_ (.A1(_1103_),
    .A2(\u1.ordering_complete[12] ),
    .B(_1105_),
    .C(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1483_ (.A1(_1099_),
    .A2(_1102_),
    .A3(_1107_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1484_ (.I(\u1.ordering_timer[9] ),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1485_ (.I(\u1.ordering_complete[9] ),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1486_ (.I(\u1.ordering_timer[8] ),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1487_ (.I(\u1.ordering_complete[8] ),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1488_ (.I(\u1.ordering_complete[10] ),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1489_ (.A1(\u1.ordering_timer[11] ),
    .A2(_1104_),
    .B1(\u1.ordering_timer[10] ),
    .B2(_1113_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1490_ (.A1(_1109_),
    .A2(_1110_),
    .B1(_1111_),
    .B2(_1112_),
    .C(_1114_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1491_ (.I(\u1.ordering_timer[10] ),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1492_ (.A1(_1116_),
    .A2(\u1.ordering_complete[10] ),
    .B1(_1109_),
    .B2(\u1.ordering_complete[9] ),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1493_ (.A1(_1111_),
    .A2(_1112_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1494_ (.A1(_1117_),
    .A2(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1495_ (.A1(_1108_),
    .A2(_1115_),
    .A3(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1496_ (.I(\u1.ordering_timer[5] ),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1497_ (.I(\u1.ordering_timer[4] ),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1498_ (.A1(_1121_),
    .A2(\u1.ordering_complete[5] ),
    .B1(_1122_),
    .B2(\u1.ordering_complete[4] ),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1499_ (.I(\u1.ordering_timer[7] ),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1500_ (.I(\u1.ordering_timer[6] ),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1501_ (.A1(_1124_),
    .A2(\u1.ordering_complete[7] ),
    .B1(_1125_),
    .B2(\u1.ordering_complete[6] ),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1502_ (.A1(_1123_),
    .A2(_1126_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1503_ (.I(\u1.ordering_timer[3] ),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1504_ (.A1(_1124_),
    .A2(\u1.ordering_complete[7] ),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1505_ (.A1(_1128_),
    .A2(\u1.ordering_complete[3] ),
    .B1(_1122_),
    .B2(\u1.ordering_complete[4] ),
    .C(_1129_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1506_ (.A1(_1125_),
    .A2(\u1.ordering_complete[6] ),
    .B1(_1121_),
    .B2(\u1.ordering_complete[5] ),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1507_ (.A1(_1127_),
    .A2(_1130_),
    .A3(_1131_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1508_ (.I(\u1.ordering_complete[0] ),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1509_ (.I(\u1.ordering_complete[1] ),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1510_ (.A1(\u1.ordering_timer[0] ),
    .A2(_1133_),
    .B1(\u1.ordering_timer[1] ),
    .B2(_1134_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1511_ (.I(\u1.ordering_timer[2] ),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1512_ (.A1(_1128_),
    .A2(\u1.ordering_complete[3] ),
    .B1(_1136_),
    .B2(\u1.ordering_complete[2] ),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1513_ (.I(\u1.ordering_timer[0] ),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1514_ (.I(_1138_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1515_ (.A1(\u1.ordering_timer[1] ),
    .A2(_1134_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1516_ (.A1(_1136_),
    .A2(\u1.ordering_complete[2] ),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1517_ (.A1(_1139_),
    .A2(\u1.ordering_complete[0] ),
    .B(_1140_),
    .C(_1141_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1518_ (.A1(_1132_),
    .A2(_1135_),
    .A3(_1137_),
    .A4(_1142_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1519_ (.A1(_1070_),
    .A2(_1095_),
    .A3(_1120_),
    .A4(_1143_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1520_ (.I(_1144_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1521_ (.A1(\u0.run_state[6] ),
    .A2(_1045_),
    .B1(_1145_),
    .B2(\u0.run_state[3] ),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1522_ (.A1(_1043_),
    .A2(_1146_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1523_ (.A1(\control_trigger_sync[0] ),
    .A2(control_trigger),
    .A3(\control_trigger_sync[1] ),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1524_ (.A1(\u0.cmd[28] ),
    .A2(\u0.run_state[2] ),
    .B1(_1147_),
    .B2(\u0.run_state[5] ),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1525_ (.A1(_1043_),
    .A2(_1148_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1526_ (.I(\u0.cmd[27] ),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1527_ (.A1(\u0.run_state[5] ),
    .A2(_1044_),
    .B(\u0.run_state[1] ),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1528_ (.A1(_1149_),
    .A2(_1150_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1529_ (.A1(\u0.run_state[4] ),
    .A2(_1151_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1530_ (.A1(_1043_),
    .A2(_1152_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1531_ (.I(\u0.cmd[29] ),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1532_ (.I(\u0.run_state[0] ),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1533_ (.A1(_1040_),
    .A2(\u0.cmd[30] ),
    .A3(_1042_),
    .Z(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1534_ (.A1(_1153_),
    .A2(_1154_),
    .B(_1155_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1535_ (.I(\u0.u11.impulse_gen[0] ),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1536_ (.A1(_1156_),
    .A2(\u0.u11.impulse_gen[1] ),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1537_ (.I(_1157_),
    .Z(\u0.latch_cmd ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1538_ (.A1(\u0.run_state[3] ),
    .A2(\u0.run_state[4] ),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1539_ (.I(_1158_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1540_ (.I(\u0.run_state[6] ),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1541_ (.I(\u0.cmd[27] ),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1542_ (.A1(_1159_),
    .A2(_1045_),
    .B1(_1150_),
    .B2(_1160_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1543_ (.A1(\u0.run_state[3] ),
    .A2(_1144_),
    .B(_1161_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1544_ (.A1(_1043_),
    .A2(_1162_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1545_ (.I(\u1.timer[25] ),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1546_ (.I(_1163_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1547_ (.I(\u1.timer[24] ),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1548_ (.I(_1165_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1549_ (.I(\u1.timer[30] ),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1550_ (.I(\u1.timer[29] ),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1551_ (.A1(\u1.ccr1[30] ),
    .A2(_1167_),
    .B1(\u1.ccr1[29] ),
    .B2(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1552_ (.A1(\u1.ccr1[25] ),
    .A2(_1164_),
    .B1(\u1.ccr1[24] ),
    .B2(_1166_),
    .C(_1169_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1553_ (.I(\u1.timer[31] ),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1554_ (.A1(\u1.ccr1[31] ),
    .A2(_1171_),
    .B1(\u1.ccr1[30] ),
    .B2(_1167_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1555_ (.I(\u1.timer[28] ),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1556_ (.A1(\u1.ccr1[29] ),
    .A2(_1168_),
    .B1(\u1.ccr1[28] ),
    .B2(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1557_ (.A1(_1172_),
    .A2(_1174_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1558_ (.I(\u1.ccr1[27] ),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1559_ (.I(\u1.timer[27] ),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1560_ (.I(\u1.ccr1[26] ),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1561_ (.A1(_1176_),
    .A2(\u1.timer[27] ),
    .B1(_1178_),
    .B2(\u1.timer[26] ),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1562_ (.I(\u1.timer[26] ),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1563_ (.A1(\u1.ccr1[26] ),
    .A2(_1180_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1564_ (.A1(_1176_),
    .A2(_1177_),
    .B(_1179_),
    .C(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1565_ (.A1(\u1.ccr1[25] ),
    .A2(_1163_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1566_ (.A1(\u1.ccr1[28] ),
    .A2(_1173_),
    .B1(\u1.ccr1[24] ),
    .B2(_1165_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1567_ (.A1(\u1.ccr1[31] ),
    .A2(_1171_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1568_ (.A1(_1183_),
    .A2(_1184_),
    .A3(_1185_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1569_ (.A1(_1170_),
    .A2(_1175_),
    .A3(_1182_),
    .A4(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1570_ (.I(\u1.timer[6] ),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1571_ (.I(_1188_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1572_ (.I(\u1.timer[5] ),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1573_ (.I(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1574_ (.A1(\u1.ccr1[6] ),
    .A2(_1189_),
    .B1(\u1.ccr1[5] ),
    .B2(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1575_ (.I(\u1.timer[7] ),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1576_ (.I(\u1.timer[4] ),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1577_ (.A1(\u1.ccr1[7] ),
    .A2(_1193_),
    .B1(\u1.ccr1[4] ),
    .B2(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1578_ (.I(\u1.ccr1[5] ),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1579_ (.I(\u1.ccr1[4] ),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1580_ (.A1(_1196_),
    .A2(_1190_),
    .B1(_1197_),
    .B2(\u1.timer[4] ),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1581_ (.I(\u1.ccr1[7] ),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1582_ (.I(\u1.ccr1[6] ),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1583_ (.A1(_1199_),
    .A2(\u1.timer[7] ),
    .B1(_1200_),
    .B2(_1188_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1584_ (.A1(_1192_),
    .A2(_1195_),
    .A3(_1198_),
    .A4(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1585_ (.I(\u1.timer[2] ),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1586_ (.I(_1203_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1587_ (.A1(\u1.ccr1[2] ),
    .A2(_1204_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1588_ (.I(\u1.timer[0] ),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1589_ (.I(_1206_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1590_ (.I(\u1.timer[1] ),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1591_ (.I(_1208_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1592_ (.A1(_1207_),
    .A2(\u1.ccr1[0] ),
    .B1(\u1.ccr1[1] ),
    .B2(_1209_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1593_ (.A1(_1205_),
    .A2(_1210_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1594_ (.I(\u0.timer_enable ),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1595_ (.I(\u1.ccr1[3] ),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1596_ (.I(\u1.timer[3] ),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1597_ (.I(\u1.ccr1[2] ),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1598_ (.A1(_1213_),
    .A2(_1214_),
    .B1(_1215_),
    .B2(_1203_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1599_ (.A1(_1207_),
    .A2(\u1.ccr1[0] ),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1600_ (.A1(\u1.ccr1[1] ),
    .A2(_1209_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1601_ (.A1(_1213_),
    .A2(\u1.timer[3] ),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1602_ (.A1(_1218_),
    .A2(_1219_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1603_ (.A1(_1212_),
    .A2(_1216_),
    .A3(_1217_),
    .A4(_1220_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1604_ (.A1(_1202_),
    .A2(_1211_),
    .A3(_1221_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1605_ (.I(\u1.timer[20] ),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1606_ (.I(_1223_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1607_ (.I(\u1.ccr1[23] ),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1608_ (.I(\u1.ccr1[22] ),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1609_ (.A1(_1225_),
    .A2(\u1.timer[23] ),
    .B1(_1226_),
    .B2(\u1.timer[22] ),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1610_ (.I(\u1.timer[23] ),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1611_ (.I(\u1.timer[22] ),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1612_ (.I(\u1.timer[21] ),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _1613_ (.A1(\u1.ccr1[23] ),
    .A2(_1228_),
    .B1(\u1.ccr1[22] ),
    .B2(_1229_),
    .C1(\u1.ccr1[21] ),
    .C2(_1230_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1614_ (.A1(_1227_),
    .A2(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1615_ (.I(_1230_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1616_ (.A1(\u1.ccr1[21] ),
    .A2(_1233_),
    .B1(\u1.ccr1[20] ),
    .B2(_1223_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1617_ (.A1(\u1.ccr1[20] ),
    .A2(_1224_),
    .B(_1232_),
    .C(_1234_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1618_ (.I(\u1.timer[17] ),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1619_ (.I(\u1.timer[16] ),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1620_ (.A1(\u1.ccr1[17] ),
    .A2(_1236_),
    .B1(\u1.ccr1[16] ),
    .B2(_1237_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1621_ (.A1(\u1.ccr1[19] ),
    .A2(\u1.timer[19] ),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1622_ (.A1(\u1.ccr1[18] ),
    .A2(\u1.timer[18] ),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1623_ (.A1(_1239_),
    .A2(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1624_ (.A1(\u1.ccr1[17] ),
    .A2(_1236_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1625_ (.A1(\u1.ccr1[16] ),
    .A2(_1237_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1626_ (.A1(_1241_),
    .A2(_1242_),
    .A3(_1243_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1627_ (.A1(_1238_),
    .A2(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1628_ (.A1(_1235_),
    .A2(_1245_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1629_ (.I(\u1.ccr1[9] ),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1630_ (.I(\u1.timer[9] ),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1631_ (.I(\u1.ccr1[8] ),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1632_ (.I(\u1.timer[8] ),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1633_ (.A1(_1247_),
    .A2(_1248_),
    .B1(_1249_),
    .B2(_1250_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1634_ (.I(\u1.ccr1[15] ),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1635_ (.I(\u1.ccr1[14] ),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1636_ (.I(\u1.timer[14] ),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1637_ (.A1(_1252_),
    .A2(\u1.timer[15] ),
    .B1(_1253_),
    .B2(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1638_ (.I(\u1.timer[15] ),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1639_ (.I(\u1.timer[14] ),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1640_ (.I(\u1.timer[13] ),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1641_ (.A1(\u1.ccr1[15] ),
    .A2(_1256_),
    .B1(\u1.ccr1[14] ),
    .B2(_1257_),
    .C1(\u1.ccr1[13] ),
    .C2(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1642_ (.A1(_1255_),
    .A2(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1643_ (.I(\u1.ccr1[12] ),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1644_ (.I(\u1.timer[12] ),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1645_ (.I(\u1.ccr1[13] ),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1646_ (.A1(_1263_),
    .A2(\u1.timer[13] ),
    .B1(_1261_),
    .B2(\u1.timer[12] ),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1647_ (.A1(_1261_),
    .A2(_1262_),
    .B(_1264_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1648_ (.A1(_1260_),
    .A2(_1265_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1649_ (.I(\u1.timer[8] ),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1650_ (.I(\u1.timer[10] ),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1651_ (.I(\u1.timer[11] ),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1652_ (.A1(\u1.ccr1[11] ),
    .A2(_1269_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1653_ (.I(\u1.ccr1[11] ),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1654_ (.I(\u1.timer[11] ),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1655_ (.A1(_1271_),
    .A2(_1272_),
    .B1(\u1.ccr1[10] ),
    .B2(_1268_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1656_ (.A1(\u1.ccr1[10] ),
    .A2(_1268_),
    .B(_1270_),
    .C(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1657_ (.A1(_1247_),
    .A2(_1248_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1658_ (.A1(\u1.ccr1[8] ),
    .A2(_1267_),
    .B(_1274_),
    .C(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1659_ (.A1(_1251_),
    .A2(_1266_),
    .A3(_1276_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1660_ (.A1(_1246_),
    .A2(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1661_ (.A1(_1187_),
    .A2(_1222_),
    .A3(_1278_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1662_ (.I(_1279_),
    .ZN(\u1.ccr1_flag ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1663_ (.I(_1188_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1664_ (.I(\u1.ccr0[6] ),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1665_ (.I(\u1.ccr0[5] ),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1666_ (.I(_1190_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1667_ (.A1(_1280_),
    .A2(_1281_),
    .B1(_1282_),
    .B2(_1283_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1668_ (.A1(_1193_),
    .A2(\u1.ccr0[7] ),
    .B1(\u1.ccr0[4] ),
    .B2(_1194_),
    .C(_1284_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1669_ (.I(\u1.ccr0[4] ),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1670_ (.I(\u1.timer[4] ),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1671_ (.A1(_1283_),
    .A2(_1282_),
    .B1(_1286_),
    .B2(_1287_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1672_ (.I(\u1.timer[7] ),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1673_ (.I(\u1.ccr0[7] ),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1674_ (.A1(_1289_),
    .A2(_1290_),
    .B1(_1281_),
    .B2(_1280_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1675_ (.A1(_1285_),
    .A2(_1288_),
    .A3(_1291_),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1676_ (.I(\u1.timer[9] ),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1677_ (.A1(_1269_),
    .A2(\u1.ccr0[11] ),
    .B1(\u1.ccr0[10] ),
    .B2(_1268_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1678_ (.I(\u1.timer[10] ),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1679_ (.I(\u1.ccr0[10] ),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1680_ (.A1(_1269_),
    .A2(\u1.ccr0[11] ),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1681_ (.A1(_1295_),
    .A2(_1296_),
    .B(_1297_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1682_ (.A1(_1293_),
    .A2(\u1.ccr0[9] ),
    .B(_1294_),
    .C(_1298_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1683_ (.I(\u1.timer[13] ),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1684_ (.I(\u1.ccr0[13] ),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1685_ (.A1(_1300_),
    .A2(_1301_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1686_ (.I(\u1.timer[15] ),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1687_ (.I(\u1.ccr0[15] ),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1688_ (.I(\u1.ccr0[14] ),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1689_ (.A1(_1303_),
    .A2(_1304_),
    .B1(_1305_),
    .B2(_1254_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1690_ (.A1(_1256_),
    .A2(\u1.ccr0[15] ),
    .B1(\u1.ccr0[14] ),
    .B2(_1257_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1691_ (.A1(_1306_),
    .A2(_1307_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1692_ (.A1(_1293_),
    .A2(\u1.ccr0[9] ),
    .B1(\u1.ccr0[8] ),
    .B2(_1267_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1693_ (.I(\u1.ccr0[12] ),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1694_ (.I(_1262_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1695_ (.A1(_1300_),
    .A2(_1301_),
    .B1(_1310_),
    .B2(_1311_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1696_ (.A1(_1262_),
    .A2(_1310_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1697_ (.A1(_1267_),
    .A2(\u1.ccr0[8] ),
    .B(_1313_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1698_ (.A1(_1312_),
    .A2(_1314_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1699_ (.A1(_1302_),
    .A2(_1308_),
    .A3(_1309_),
    .A4(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1700_ (.A1(_1299_),
    .A2(_1316_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1701_ (.I(\u1.timer[19] ),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1702_ (.I(\u1.ccr0[19] ),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1703_ (.I(\u1.ccr0[18] ),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1704_ (.I(\u1.timer[18] ),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1705_ (.I(_1321_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1706_ (.A1(_1318_),
    .A2(_1319_),
    .B1(_1320_),
    .B2(_1322_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1707_ (.A1(_1321_),
    .A2(_1320_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1708_ (.A1(_1318_),
    .A2(_1319_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1709_ (.A1(_1324_),
    .A2(_1325_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1710_ (.I(\u1.timer[23] ),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1711_ (.I(\u1.ccr0[23] ),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1712_ (.I(\u1.ccr0[22] ),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1713_ (.A1(_1327_),
    .A2(_1328_),
    .B1(_1329_),
    .B2(\u1.timer[22] ),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1714_ (.A1(_1327_),
    .A2(_1328_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1715_ (.A1(_1229_),
    .A2(\u1.ccr0[22] ),
    .B(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1716_ (.A1(_1330_),
    .A2(_1332_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1717_ (.A1(_1236_),
    .A2(\u1.ccr0[17] ),
    .B1(\u1.ccr0[16] ),
    .B2(_1237_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1718_ (.A1(_1233_),
    .A2(\u1.ccr0[21] ),
    .B1(\u1.ccr0[20] ),
    .B2(_1224_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1719_ (.A1(_1236_),
    .A2(\u1.ccr0[17] ),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1720_ (.A1(_1233_),
    .A2(\u1.ccr0[21] ),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1721_ (.A1(_1224_),
    .A2(\u1.ccr0[20] ),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1722_ (.A1(_1237_),
    .A2(\u1.ccr0[16] ),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1723_ (.A1(_1336_),
    .A2(_1337_),
    .A3(_1338_),
    .A4(_1339_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1724_ (.A1(_1333_),
    .A2(_1334_),
    .A3(_1335_),
    .A4(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1725_ (.A1(_1323_),
    .A2(_1326_),
    .A3(_1341_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1726_ (.I(\u1.ccr0[27] ),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1727_ (.I(\u1.ccr0[26] ),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1728_ (.I(\u1.timer[26] ),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1729_ (.A1(_1177_),
    .A2(_1343_),
    .B1(_1344_),
    .B2(_1345_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1730_ (.A1(_1164_),
    .A2(\u1.ccr0[25] ),
    .B1(\u1.ccr0[24] ),
    .B2(_1166_),
    .C(_1346_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1731_ (.A1(_1180_),
    .A2(\u1.ccr0[26] ),
    .B1(\u1.ccr0[25] ),
    .B2(_1164_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1732_ (.I(_1177_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1733_ (.A1(_1173_),
    .A2(\u1.ccr0[28] ),
    .B1(\u1.ccr0[27] ),
    .B2(_1349_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1734_ (.I(\u1.timer[31] ),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1735_ (.I(\u1.ccr0[31] ),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1736_ (.I(\u1.ccr0[30] ),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1737_ (.A1(_1351_),
    .A2(_1352_),
    .B1(_1353_),
    .B2(\u1.timer[30] ),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1738_ (.A1(_1171_),
    .A2(\u1.ccr0[31] ),
    .B1(\u1.ccr0[24] ),
    .B2(_1166_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1739_ (.A1(_1348_),
    .A2(_1350_),
    .A3(_1354_),
    .A4(_1355_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1740_ (.I(\u1.ccr0[29] ),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1741_ (.I(\u1.ccr0[28] ),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1742_ (.A1(\u1.timer[29] ),
    .A2(_1357_),
    .B1(_1358_),
    .B2(\u1.timer[28] ),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1743_ (.A1(_1167_),
    .A2(\u1.ccr0[30] ),
    .B1(\u1.ccr0[29] ),
    .B2(_1168_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1744_ (.A1(_1359_),
    .A2(_1360_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1745_ (.A1(_1347_),
    .A2(_1356_),
    .A3(_1361_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1746_ (.I(_1209_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1747_ (.I(_1207_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1748_ (.A1(_1363_),
    .A2(\u1.ccr0[1] ),
    .B1(\u1.ccr0[0] ),
    .B2(_1364_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1749_ (.A1(_1363_),
    .A2(\u1.ccr0[1] ),
    .B(_1365_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1750_ (.I(_1214_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1751_ (.A1(_1367_),
    .A2(\u1.ccr0[3] ),
    .B1(\u1.ccr0[2] ),
    .B2(_1204_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1752_ (.A1(_1367_),
    .A2(\u1.ccr0[3] ),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1753_ (.A1(_1204_),
    .A2(\u1.ccr0[2] ),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1754_ (.A1(_1364_),
    .A2(\u1.ccr0[0] ),
    .B(_1369_),
    .C(_1370_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1755_ (.A1(_1366_),
    .A2(_1368_),
    .A3(_1371_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1756_ (.A1(_1362_),
    .A2(_1372_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1757_ (.A1(_1317_),
    .A2(_1342_),
    .A3(_1373_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1758_ (.A1(_1299_),
    .A2(_1316_),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1759_ (.A1(_1363_),
    .A2(\u1.ccr0[1] ),
    .B(_1366_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1760_ (.A1(_1370_),
    .A2(_1376_),
    .B(_1368_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1761_ (.A1(_1292_),
    .A2(_1369_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1762_ (.A1(_1284_),
    .A2(_1288_),
    .B(_1291_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1763_ (.A1(_1289_),
    .A2(_1290_),
    .B(_1379_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1764_ (.A1(_1377_),
    .A2(_1378_),
    .B(_1380_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1765_ (.A1(_1294_),
    .A2(_1297_),
    .B1(_1299_),
    .B2(_1309_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1766_ (.A1(_1313_),
    .A2(_1382_),
    .B(_1312_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1767_ (.A1(_1302_),
    .A2(_1308_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1768_ (.A1(_1256_),
    .A2(\u1.ccr0[15] ),
    .B(_1306_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1769_ (.A1(_1375_),
    .A2(_1381_),
    .B1(_1383_),
    .B2(_1384_),
    .C(_1385_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1770_ (.A1(_1323_),
    .A2(_1326_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1771_ (.A1(_1336_),
    .A2(_1334_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1772_ (.A1(_1323_),
    .A2(_1325_),
    .B1(_1387_),
    .B2(_1388_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1773_ (.A1(_1338_),
    .A2(_1389_),
    .B(_1335_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1774_ (.A1(_1333_),
    .A2(_1390_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1775_ (.A1(_1337_),
    .A2(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1776_ (.A1(_1330_),
    .A2(_1331_),
    .B1(_1342_),
    .B2(_1386_),
    .C(_1392_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1777_ (.I(_1177_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1778_ (.A1(_1394_),
    .A2(_1343_),
    .B1(_1344_),
    .B2(_1345_),
    .C(_1348_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1779_ (.A1(_1350_),
    .A2(_1347_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1780_ (.A1(_1395_),
    .A2(_1396_),
    .B(_1359_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1781_ (.A1(_1360_),
    .A2(_1397_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1782_ (.A1(_1171_),
    .A2(\u1.ccr0[31] ),
    .B1(_1354_),
    .B2(_1398_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1783_ (.A1(_1362_),
    .A2(_1393_),
    .B(_1399_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1784_ (.A1(_1292_),
    .A2(_1374_),
    .B(_1400_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1785_ (.I(\u0.timer_enable ),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1786_ (.A1(_1402_),
    .A2(_1144_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1787_ (.I(_1311_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1788_ (.A1(_1256_),
    .A2(_1257_),
    .A3(_1258_),
    .A4(_1404_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1789_ (.A1(_1289_),
    .A2(_1280_),
    .A3(_1283_),
    .A4(_1287_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1790_ (.A1(_1206_),
    .A2(_1208_),
    .A3(_1214_),
    .A4(_1203_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1791_ (.A1(_1272_),
    .A2(_1295_),
    .A3(_1248_),
    .A4(_1250_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1792_ (.A1(_1406_),
    .A2(_1407_),
    .A3(_1408_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1793_ (.I(_1345_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1794_ (.I(\u1.timer[25] ),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1795_ (.A1(_1394_),
    .A2(_1410_),
    .A3(_1411_),
    .A4(\u1.timer[24] ),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1796_ (.I(\u1.timer[28] ),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1797_ (.A1(_1351_),
    .A2(\u1.timer[30] ),
    .A3(\u1.timer[29] ),
    .A4(_1413_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1798_ (.A1(_1412_),
    .A2(_1414_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1799_ (.I(_1318_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1800_ (.I(\u1.timer[17] ),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1801_ (.I(\u1.timer[16] ),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1802_ (.A1(_0281_),
    .A2(_1322_),
    .A3(_0282_),
    .A4(_0283_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1803_ (.I(_1327_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1804_ (.I(\u1.timer[22] ),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1805_ (.A1(_0285_),
    .A2(_0286_),
    .A3(\u1.timer[21] ),
    .A4(\u1.timer[20] ),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1806_ (.A1(_0284_),
    .A2(_0287_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1807_ (.A1(_1405_),
    .A2(_1409_),
    .A3(_0280_),
    .A4(_0288_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1808_ (.A1(_1401_),
    .A2(_1403_),
    .A3(_0289_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1809_ (.I0(net16),
    .I1(net3),
    .S(net34),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1810_ (.I(_0290_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1811_ (.I0(net17),
    .I1(net2),
    .S(net35),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1812_ (.I(_0291_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1813_ (.I0(net18),
    .I1(net1),
    .S(net36),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1814_ (.I(_0292_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1815_ (.A1(net19),
    .A2(net37),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1816_ (.A1(net37),
    .A2(_1144_),
    .B(_0293_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1817_ (.A1(\u0.cmd[29] ),
    .A2(\u0.run_state[0] ),
    .A3(_1155_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1818_ (.I(_0294_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1819_ (.I(\u0.cmd[30] ),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1820_ (.A1(_1040_),
    .A2(_0295_),
    .A3(\u0.update_cmd ),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1821_ (.A1(\u0.cmd[28] ),
    .A2(\u0.cmd[29] ),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1822_ (.A1(_0295_),
    .A2(\u0.update_cmd ),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1823_ (.A1(\u0.cmd[31] ),
    .A2(\u0.cmd[26] ),
    .A3(\u0.cmd[27] ),
    .A4(_0297_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1824_ (.A1(_0296_),
    .A2(_0298_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1825_ (.I(\u0.cmd[26] ),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1826_ (.A1(\u0.cmd[31] ),
    .A2(_0297_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1827_ (.A1(_0299_),
    .A2(_1149_),
    .A3(_0300_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1828_ (.A1(_0296_),
    .A2(_0301_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1829_ (.I(_0300_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1830_ (.A1(\u0.cmd[26] ),
    .A2(_1149_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1831_ (.A1(_0296_),
    .A2(_0302_),
    .A3(_0303_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1832_ (.A1(_0299_),
    .A2(_1160_),
    .A3(_0296_),
    .A4(_0302_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1833_ (.I(\u0.cmd[28] ),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1834_ (.A1(_0304_),
    .A2(\u0.cmd[29] ),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1835_ (.A1(_0298_),
    .A2(_0305_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1836_ (.A1(_0301_),
    .A2(_0305_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1837_ (.A1(_0302_),
    .A2(_0303_),
    .A3(_0305_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1838_ (.A1(_0299_),
    .A2(_1160_),
    .A3(_0302_),
    .A4(_0305_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1839_ (.A1(_0304_),
    .A2(_1153_),
    .A3(_0298_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1840_ (.A1(_0304_),
    .A2(_1153_),
    .A3(_0301_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1841_ (.A1(_0304_),
    .A2(\u0.run_state[2] ),
    .A3(_1155_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1842_ (.I(_0306_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1843_ (.I(net15),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1844_ (.A1(_0307_),
    .A2(net33),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1845_ (.I(\u1.u1.impulse_gen[1] ),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1846_ (.A1(\u1.u1.impulse_gen[0] ),
    .A2(_0308_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1847_ (.I(\u1.col_limit[6] ),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1848_ (.I(\u1.col_sel[5] ),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1849_ (.A1(_0311_),
    .A2(\u1.col_limit[5] ),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1850_ (.I(\u1.col_sel[3] ),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1851_ (.I(\u1.col_sel[4] ),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1852_ (.A1(_0313_),
    .A2(\u1.col_limit[3] ),
    .B1(_0314_),
    .B2(\u1.col_limit[4] ),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1853_ (.I(\u1.col_sel[2] ),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1854_ (.I(\u1.col_sel[1] ),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1855_ (.I(\u1.col_limit[1] ),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1856_ (.I(\u1.col_limit[2] ),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1857_ (.A1(_0317_),
    .A2(_0318_),
    .B1(\u1.col_sel[2] ),
    .B2(_0319_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1858_ (.I(\u1.col_limit[0] ),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1859_ (.A1(\u1.col_sel[0] ),
    .A2(_0321_),
    .B1(\u1.col_sel[1] ),
    .B2(_0318_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1860_ (.A1(_0313_),
    .A2(\u1.col_limit[3] ),
    .B1(_0316_),
    .B2(\u1.col_limit[2] ),
    .C1(_0320_),
    .C2(_0322_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1861_ (.A1(_0311_),
    .A2(\u1.col_limit[5] ),
    .B1(_0314_),
    .B2(\u1.col_limit[4] ),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1862_ (.A1(_0315_),
    .A2(_0323_),
    .B(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1863_ (.A1(\u1.col_sel[6] ),
    .A2(\u1.col_limit[6] ),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1864_ (.A1(_0312_),
    .A2(_0325_),
    .B(_0326_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1865_ (.A1(\u1.col_sel[6] ),
    .A2(_0310_),
    .B(_0327_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1866_ (.I(_1402_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1867_ (.A1(_0309_),
    .A2(_0328_),
    .B(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1868_ (.I(_0330_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1869_ (.A1(_1212_),
    .A2(_0309_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1870_ (.A1(\u1.col_sel[0] ),
    .A2(_0332_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1871_ (.A1(\u1.col_sel[0] ),
    .A2(_0332_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1872_ (.A1(_0331_),
    .A2(_0333_),
    .A3(_0334_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1873_ (.A1(_0317_),
    .A2(_0333_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1874_ (.A1(_0331_),
    .A2(_0335_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1875_ (.A1(_0317_),
    .A2(\u1.col_sel[2] ),
    .A3(_0333_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1876_ (.A1(_0317_),
    .A2(_0333_),
    .B(\u1.col_sel[2] ),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1877_ (.A1(_0330_),
    .A2(_0336_),
    .A3(_0337_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1878_ (.A1(\u1.col_sel[3] ),
    .A2(_0336_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1879_ (.A1(\u1.col_sel[3] ),
    .A2(_0336_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1880_ (.A1(_0330_),
    .A2(_0338_),
    .A3(_0339_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1881_ (.A1(\u1.col_sel[4] ),
    .A2(_0338_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1882_ (.A1(\u1.col_sel[4] ),
    .A2(_0338_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1883_ (.A1(_0330_),
    .A2(_0340_),
    .A3(_0341_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1884_ (.A1(_0311_),
    .A2(_0340_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1885_ (.A1(_0331_),
    .A2(_0342_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1886_ (.A1(\u1.col_sel[5] ),
    .A2(_0340_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1887_ (.A1(\u1.col_sel[6] ),
    .A2(_0343_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1888_ (.A1(_0331_),
    .A2(_0344_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1889_ (.I(\u0.cmd[0] ),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1890_ (.I(\u0.cmd[16] ),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1891_ (.I(\u0.cmd[17] ),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1892_ (.I(_0347_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1893_ (.I(\u0.cmd[19] ),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1894_ (.A1(\u0.write_config_n ),
    .A2(\u0.cmd[18] ),
    .A3(\u0.cmd[21] ),
    .A4(\u0.cmd[20] ),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1895_ (.A1(_0349_),
    .A2(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1896_ (.A1(_0346_),
    .A2(_0348_),
    .A3(_0351_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1897_ (.I(_0352_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1898_ (.I(_0353_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1899_ (.I0(\u1.ccr0[16] ),
    .I1(_0345_),
    .S(_0354_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1900_ (.I(_0355_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1901_ (.I(\u0.cmd[1] ),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1902_ (.I0(\u1.ccr0[17] ),
    .I1(_0356_),
    .S(_0354_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1903_ (.I(_0357_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1904_ (.I(_0352_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1905_ (.I(_0358_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1906_ (.I(\u0.cmd[2] ),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1907_ (.I(_0353_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1908_ (.A1(_0360_),
    .A2(_0361_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1909_ (.A1(_1320_),
    .A2(_0359_),
    .B(_0362_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1910_ (.I(\u0.cmd[3] ),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1911_ (.A1(_0363_),
    .A2(_0361_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1912_ (.A1(_1319_),
    .A2(_0359_),
    .B(_0364_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1913_ (.I(\u0.cmd[4] ),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1914_ (.I0(\u1.ccr0[20] ),
    .I1(_0365_),
    .S(_0354_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1915_ (.I(_0366_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1916_ (.I(\u0.cmd[5] ),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1917_ (.I0(\u1.ccr0[21] ),
    .I1(_0367_),
    .S(_0354_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1918_ (.I(_0368_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1919_ (.I(\u0.cmd[6] ),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1920_ (.I(_0353_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1921_ (.A1(_0369_),
    .A2(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1922_ (.A1(_1329_),
    .A2(_0359_),
    .B(_0371_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1923_ (.I(\u0.cmd[7] ),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1924_ (.A1(_0372_),
    .A2(_0370_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1925_ (.A1(_1328_),
    .A2(_0359_),
    .B(_0373_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1926_ (.I(\u0.cmd[8] ),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1927_ (.I0(\u1.ccr0[24] ),
    .I1(_0374_),
    .S(_0358_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1928_ (.I(_0375_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1929_ (.I(\u0.cmd[9] ),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1930_ (.I0(\u1.ccr0[25] ),
    .I1(_0376_),
    .S(_0358_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1931_ (.I(_0377_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1932_ (.I(_0358_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1933_ (.I(\u0.cmd[10] ),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1934_ (.A1(_0379_),
    .A2(_0370_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1935_ (.A1(_1344_),
    .A2(_0378_),
    .B(_0380_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1936_ (.I(\u0.cmd[11] ),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1937_ (.A1(_0381_),
    .A2(_0370_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1938_ (.A1(_1343_),
    .A2(_0378_),
    .B(_0382_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1939_ (.I(_0353_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1940_ (.A1(\u0.cmd[12] ),
    .A2(_0383_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1941_ (.A1(_1358_),
    .A2(_0378_),
    .B(_0384_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1942_ (.I(\u0.cmd[13] ),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1943_ (.A1(_0385_),
    .A2(_0383_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1944_ (.A1(_1357_),
    .A2(_0378_),
    .B(_0386_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1945_ (.I(\u0.cmd[14] ),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1946_ (.A1(_0387_),
    .A2(_0383_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1947_ (.A1(_1353_),
    .A2(_0361_),
    .B(_0388_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1948_ (.I(\u0.cmd[15] ),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1949_ (.A1(_0389_),
    .A2(_0383_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1950_ (.A1(_1352_),
    .A2(_0361_),
    .B(_0390_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1951_ (.I(\u0.cmd[17] ),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1952_ (.A1(\u0.cmd[16] ),
    .A2(_0391_),
    .A3(_0351_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1953_ (.I(_0392_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1954_ (.I(_0393_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1955_ (.I0(\u1.ccr1[0] ),
    .I1(_0345_),
    .S(_0394_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1956_ (.I(_0395_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1957_ (.I0(\u1.ccr1[1] ),
    .I1(_0356_),
    .S(_0394_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1958_ (.I(_0396_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1959_ (.I(_0393_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1960_ (.I(_0397_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1961_ (.I(\u0.cmd[2] ),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1962_ (.I(_0392_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1963_ (.A1(_0399_),
    .A2(_0400_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1964_ (.A1(_1215_),
    .A2(_0398_),
    .B(_0401_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1965_ (.I(\u0.cmd[3] ),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1966_ (.A1(_0402_),
    .A2(_0400_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1967_ (.A1(_1213_),
    .A2(_0398_),
    .B(_0403_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1968_ (.I(\u0.cmd[4] ),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1969_ (.A1(_0404_),
    .A2(_0400_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1970_ (.A1(_1197_),
    .A2(_0398_),
    .B(_0405_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1971_ (.I(\u0.cmd[5] ),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1972_ (.I(_0393_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1973_ (.A1(_0406_),
    .A2(_0407_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1974_ (.A1(_1196_),
    .A2(_0398_),
    .B(_0408_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1975_ (.I(_0397_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1976_ (.A1(_0369_),
    .A2(_0407_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1977_ (.A1(_1200_),
    .A2(_0409_),
    .B(_0410_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1978_ (.A1(_0372_),
    .A2(_0407_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1979_ (.A1(_1199_),
    .A2(_0409_),
    .B(_0411_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1980_ (.A1(\u0.cmd[8] ),
    .A2(_0407_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1981_ (.A1(_1249_),
    .A2(_0409_),
    .B(_0412_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1982_ (.I(_0393_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1983_ (.A1(\u0.cmd[9] ),
    .A2(_0413_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1984_ (.A1(_1247_),
    .A2(_0409_),
    .B(_0414_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1985_ (.I0(\u1.ccr1[10] ),
    .I1(_0379_),
    .S(_0397_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1986_ (.I(_0415_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1987_ (.I(_0397_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1988_ (.A1(_0381_),
    .A2(_0413_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1989_ (.A1(_1271_),
    .A2(_0416_),
    .B(_0417_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1990_ (.A1(\u0.cmd[12] ),
    .A2(_0413_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1991_ (.A1(_1261_),
    .A2(_0416_),
    .B(_0418_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1992_ (.A1(\u0.cmd[13] ),
    .A2(_0413_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1993_ (.A1(_1263_),
    .A2(_0416_),
    .B(_0419_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1994_ (.A1(_0387_),
    .A2(_0394_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1995_ (.A1(_1253_),
    .A2(_0416_),
    .B(_0420_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1996_ (.A1(_0389_),
    .A2(_0394_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1997_ (.A1(_1252_),
    .A2(_0400_),
    .B(_0421_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1998_ (.A1(_0346_),
    .A2(_0391_),
    .A3(_0351_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1999_ (.I(_0422_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2000_ (.I0(\u1.ccr1[16] ),
    .I1(_0345_),
    .S(_0423_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2001_ (.I(_0424_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2002_ (.I0(\u1.ccr1[17] ),
    .I1(_0356_),
    .S(_0423_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2003_ (.I(_0425_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2004_ (.I(_0422_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2005_ (.I(_0426_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2006_ (.I0(\u1.ccr1[18] ),
    .I1(_0360_),
    .S(_0427_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2007_ (.I(_0428_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2008_ (.I(\u1.ccr1[19] ),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2009_ (.I(_0426_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2010_ (.I(_0422_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2011_ (.A1(_0402_),
    .A2(_0431_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2012_ (.A1(_0429_),
    .A2(_0430_),
    .B(_0432_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2013_ (.I0(\u1.ccr1[20] ),
    .I1(_0365_),
    .S(_0427_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2014_ (.I(_0433_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2015_ (.I0(\u1.ccr1[21] ),
    .I1(_0367_),
    .S(_0427_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2016_ (.I(_0434_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2017_ (.A1(_0369_),
    .A2(_0431_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2018_ (.A1(_1226_),
    .A2(_0430_),
    .B(_0435_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2019_ (.A1(_0372_),
    .A2(_0431_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2020_ (.A1(_1225_),
    .A2(_0430_),
    .B(_0436_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2021_ (.I0(\u1.ccr1[24] ),
    .I1(_0374_),
    .S(_0427_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2022_ (.I(_0437_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2023_ (.I(_0426_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2024_ (.I0(\u1.ccr1[25] ),
    .I1(_0376_),
    .S(_0438_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2025_ (.I(_0439_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2026_ (.A1(_0379_),
    .A2(_0423_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2027_ (.A1(_1178_),
    .A2(_0430_),
    .B(_0440_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2028_ (.A1(_0381_),
    .A2(_0423_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2029_ (.A1(_1176_),
    .A2(_0431_),
    .B(_0441_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2030_ (.I(\u0.cmd[12] ),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2031_ (.I0(\u1.ccr1[28] ),
    .I1(_0442_),
    .S(_0438_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2032_ (.I(_0443_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2033_ (.I0(\u1.ccr1[29] ),
    .I1(_0385_),
    .S(_0438_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2034_ (.I(_0444_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2035_ (.I0(\u1.ccr1[30] ),
    .I1(_0387_),
    .S(_0438_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2036_ (.I(_0445_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2037_ (.I0(\u1.ccr1[31] ),
    .I1(_0389_),
    .S(_0426_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2038_ (.I(_0446_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2039_ (.I(\u0.cmd[16] ),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2040_ (.A1(_0447_),
    .A2(_0347_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2041_ (.A1(\u0.cmd[18] ),
    .A2(_0349_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2042_ (.A1(\u0.write_config_n ),
    .A2(\u0.cmd[21] ),
    .A3(\u0.cmd[20] ),
    .A4(_0449_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2043_ (.A1(_0448_),
    .A2(_0450_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2044_ (.I(_0451_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2045_ (.I(_0452_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2046_ (.I(\u0.cmd[0] ),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2047_ (.I(_0451_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2048_ (.A1(_0454_),
    .A2(_0455_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2049_ (.A1(_1133_),
    .A2(_0453_),
    .B(_0456_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2050_ (.I(\u0.cmd[1] ),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2051_ (.A1(_0457_),
    .A2(_0455_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2052_ (.A1(_1134_),
    .A2(_0453_),
    .B(_0458_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2053_ (.I(_0399_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2054_ (.I(_0452_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2055_ (.I0(_0459_),
    .I1(\u1.ordering_complete[2] ),
    .S(_0460_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2056_ (.I(_0461_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2057_ (.I(_0402_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2058_ (.I0(_0462_),
    .I1(\u1.ordering_complete[3] ),
    .S(_0460_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2059_ (.I(_0463_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2060_ (.I(_0404_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2061_ (.I0(_0464_),
    .I1(\u1.ordering_complete[4] ),
    .S(_0460_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2062_ (.I(_0465_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2063_ (.I(_0406_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2064_ (.I0(_0466_),
    .I1(\u1.ordering_complete[5] ),
    .S(_0460_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2065_ (.I(_0467_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2066_ (.I(\u0.cmd[6] ),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2067_ (.I(_0468_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2068_ (.I(_0451_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2069_ (.I0(_0469_),
    .I1(\u1.ordering_complete[6] ),
    .S(_0470_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2070_ (.I(_0471_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2071_ (.I(\u0.cmd[7] ),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2072_ (.I0(_0472_),
    .I1(\u1.ordering_complete[7] ),
    .S(_0470_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2073_ (.I(_0473_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2074_ (.I(\u0.cmd[8] ),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2075_ (.I0(_0474_),
    .I1(_1112_),
    .S(_0470_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2076_ (.I(_0475_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2077_ (.I(\u0.cmd[9] ),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2078_ (.I0(_0476_),
    .I1(_1110_),
    .S(_0470_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2079_ (.I(_0477_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2080_ (.I(_0451_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2081_ (.A1(\u0.cmd[10] ),
    .A2(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2082_ (.A1(_1113_),
    .A2(_0453_),
    .B(_0479_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2083_ (.A1(\u0.cmd[11] ),
    .A2(_0478_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2084_ (.A1(_1104_),
    .A2(_0453_),
    .B(_0480_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2085_ (.I0(_0442_),
    .I1(\u1.ordering_complete[12] ),
    .S(_0452_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2086_ (.I(_0481_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2087_ (.I0(_0385_),
    .I1(\u1.ordering_complete[13] ),
    .S(_0452_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2088_ (.I(_0482_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2089_ (.A1(\u0.cmd[14] ),
    .A2(_0478_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2090_ (.A1(_1098_),
    .A2(_0455_),
    .B(_0483_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2091_ (.A1(\u0.cmd[15] ),
    .A2(_0478_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2092_ (.A1(_1097_),
    .A2(_0455_),
    .B(_0484_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2093_ (.A1(_0346_),
    .A2(_0347_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2094_ (.A1(_0485_),
    .A2(_0450_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2095_ (.I(_0486_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2096_ (.I(_0487_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2097_ (.I(_0488_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2098_ (.I(_0487_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2099_ (.A1(_0454_),
    .A2(_0490_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2100_ (.A1(_1060_),
    .A2(_0489_),
    .B(_0491_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2101_ (.A1(_0457_),
    .A2(_0490_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2102_ (.A1(_1061_),
    .A2(_0489_),
    .B(_0492_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2103_ (.I(_0487_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2104_ (.A1(_0399_),
    .A2(_0493_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2105_ (.A1(_1067_),
    .A2(_0489_),
    .B(_0494_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2106_ (.A1(_0402_),
    .A2(_0493_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2107_ (.A1(_1058_),
    .A2(_0489_),
    .B(_0495_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2108_ (.I(_0487_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2109_ (.I0(_0464_),
    .I1(\u1.ordering_complete[20] ),
    .S(_0496_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2110_ (.I(_0497_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2111_ (.I0(_0466_),
    .I1(\u1.ordering_complete[21] ),
    .S(_0496_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2112_ (.I(_0498_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2113_ (.I0(_0469_),
    .I1(\u1.ordering_complete[22] ),
    .S(_0496_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2114_ (.I(_0499_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2115_ (.I(_0488_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2116_ (.A1(\u0.cmd[7] ),
    .A2(_0493_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2117_ (.A1(_1054_),
    .A2(_0500_),
    .B(_0501_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2118_ (.I0(_0474_),
    .I1(\u1.ordering_complete[24] ),
    .S(_0496_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2119_ (.I(_0502_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2120_ (.I0(_0476_),
    .I1(\u1.ordering_complete[25] ),
    .S(_0488_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2121_ (.I(_0503_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2122_ (.I(\u1.ordering_complete[26] ),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2123_ (.A1(\u0.cmd[10] ),
    .A2(_0493_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2124_ (.A1(_0504_),
    .A2(_0500_),
    .B(_0505_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2125_ (.I(\u1.ordering_complete[27] ),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2126_ (.I(_0486_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2127_ (.A1(\u0.cmd[11] ),
    .A2(_0507_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2128_ (.A1(_0506_),
    .A2(_0500_),
    .B(_0508_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2129_ (.I0(_0442_),
    .I1(\u1.ordering_complete[28] ),
    .S(_0488_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2130_ (.I(_0509_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2131_ (.A1(\u0.cmd[13] ),
    .A2(_0507_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2132_ (.A1(_1079_),
    .A2(_0500_),
    .B(_0510_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2133_ (.A1(\u0.cmd[14] ),
    .A2(_0507_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2134_ (.A1(_1078_),
    .A2(_0490_),
    .B(_0511_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2135_ (.A1(\u0.cmd[15] ),
    .A2(_0507_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2136_ (.A1(_1073_),
    .A2(_0490_),
    .B(_0512_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2137_ (.I(_0454_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2138_ (.A1(_0346_),
    .A2(_0348_),
    .A3(_0450_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2139_ (.I(_0514_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2140_ (.I0(_0513_),
    .I1(\u1.row_limit[0] ),
    .S(_0515_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2141_ (.I(_0516_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2142_ (.I(_0457_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2143_ (.I0(_0517_),
    .I1(\u1.row_limit[1] ),
    .S(_0515_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2144_ (.I(_0518_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2145_ (.I0(_0459_),
    .I1(\u1.row_limit[2] ),
    .S(_0514_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2146_ (.I(_0519_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2147_ (.I0(_0462_),
    .I1(\u1.row_limit[3] ),
    .S(_0514_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2148_ (.I(_0520_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2149_ (.I(\u1.row_limit[4] ),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2150_ (.I(_0514_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2151_ (.A1(_0404_),
    .A2(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2152_ (.A1(_0521_),
    .A2(_0522_),
    .B(_0523_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2153_ (.I(\u1.row_limit[5] ),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2154_ (.A1(_0406_),
    .A2(_0515_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2155_ (.A1(_0524_),
    .A2(_0522_),
    .B(_0525_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2156_ (.I(\u1.row_limit[6] ),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2157_ (.A1(_0468_),
    .A2(_0515_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2158_ (.A1(_0526_),
    .A2(_0522_),
    .B(_0527_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2159_ (.A1(_0447_),
    .A2(_0348_),
    .A3(_0450_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2160_ (.I(_0528_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2161_ (.I(_0529_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2162_ (.I(_0528_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2163_ (.A1(_0454_),
    .A2(_0531_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2164_ (.A1(_0321_),
    .A2(_0530_),
    .B(_0532_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2165_ (.A1(_0457_),
    .A2(_0531_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2166_ (.A1(_0318_),
    .A2(_0530_),
    .B(_0533_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2167_ (.A1(_0399_),
    .A2(_0531_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2168_ (.A1(_0319_),
    .A2(_0530_),
    .B(_0534_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2169_ (.I0(_0462_),
    .I1(\u1.col_limit[3] ),
    .S(_0529_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2170_ (.I(_0535_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2171_ (.I0(_0464_),
    .I1(\u1.col_limit[4] ),
    .S(_0529_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2172_ (.I(_0536_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2173_ (.I0(_0466_),
    .I1(\u1.col_limit[5] ),
    .S(_0529_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2174_ (.I(_0537_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2175_ (.A1(_0468_),
    .A2(_0531_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2176_ (.A1(_0310_),
    .A2(_0530_),
    .B(_0538_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2177_ (.A1(\u0.cmd[19] ),
    .A2(_0350_),
    .A3(_0448_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2178_ (.I(_0539_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2179_ (.I0(_0513_),
    .I1(\u1.inverter_select[0] ),
    .S(_0540_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2180_ (.I(_0541_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2181_ (.I0(_0517_),
    .I1(\u1.inverter_select[1] ),
    .S(_0540_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2182_ (.I(_0542_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2183_ (.I0(_0459_),
    .I1(\u1.inverter_select[2] ),
    .S(_0540_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2184_ (.I(_0543_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2185_ (.I0(_0363_),
    .I1(\u1.inverter_select[3] ),
    .S(_0540_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2186_ (.I(_0544_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2187_ (.I(_0539_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2188_ (.I0(_0365_),
    .I1(\u1.inverter_select[4] ),
    .S(_0545_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2189_ (.I(_0546_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2190_ (.I0(_0367_),
    .I1(\u1.inverter_select[5] ),
    .S(_0545_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2191_ (.I(_0547_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2192_ (.I0(_0469_),
    .I1(\u1.inverter_select[6] ),
    .S(_0545_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2193_ (.I(_0548_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2194_ (.I0(_0472_),
    .I1(\u1.inverter_select[7] ),
    .S(_0545_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2195_ (.I(_0549_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2196_ (.I0(_0474_),
    .I1(\u1.inverter_select[8] ),
    .S(_0539_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2197_ (.I(_0550_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2198_ (.I0(_0476_),
    .I1(\u1.inverter_select[9] ),
    .S(_0539_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2199_ (.I(_0551_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2200_ (.A1(\u0.cmd[19] ),
    .A2(_0485_),
    .A3(_0350_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2201_ (.I(_0552_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2202_ (.I0(_0513_),
    .I1(\u1.row_col_select[0] ),
    .S(_0553_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2203_ (.I(_0554_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2204_ (.I0(_0517_),
    .I1(\u1.row_col_select[1] ),
    .S(_0553_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2205_ (.I(_0555_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2206_ (.I0(_0360_),
    .I1(\u1.row_col_select[2] ),
    .S(_0553_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2207_ (.I(_0556_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2208_ (.I0(_0363_),
    .I1(\u1.row_col_select[3] ),
    .S(_0553_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2209_ (.I(_0557_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2210_ (.I(_0552_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2211_ (.I0(_0365_),
    .I1(\u1.row_col_select[4] ),
    .S(_0558_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2212_ (.I(_0559_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2213_ (.I0(_0367_),
    .I1(\u1.row_col_select[5] ),
    .S(_0558_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2214_ (.I(_0560_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2215_ (.I0(_0369_),
    .I1(\u1.row_col_select[6] ),
    .S(_0558_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2216_ (.I(_0561_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2217_ (.I0(_0472_),
    .I1(\u1.row_col_select[7] ),
    .S(_0558_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2218_ (.I(_0562_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2219_ (.I0(_0374_),
    .I1(\u1.row_col_select[8] ),
    .S(_0552_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2220_ (.I(_0563_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2221_ (.I0(_0376_),
    .I1(\u1.row_col_select[9] ),
    .S(_0552_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2222_ (.I(_0564_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2223_ (.I(_1402_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2224_ (.A1(_1070_),
    .A2(_1095_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2225_ (.A1(_1135_),
    .A2(_1140_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2226_ (.A1(_1141_),
    .A2(_0567_),
    .B(_1137_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2227_ (.A1(_1123_),
    .A2(_1131_),
    .B(_1126_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2228_ (.A1(_1132_),
    .A2(_0568_),
    .B1(_0569_),
    .B2(_1129_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2229_ (.I(_1096_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2230_ (.A1(_1102_),
    .A2(_1106_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2231_ (.A1(_0571_),
    .A2(\u1.ordering_complete[15] ),
    .B1(_1099_),
    .B2(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2232_ (.A1(_1109_),
    .A2(_1110_),
    .B1(_1111_),
    .B2(\u1.ordering_complete[8] ),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2233_ (.A1(_1117_),
    .A2(_0574_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2234_ (.A1(_1114_),
    .A2(_0575_),
    .B(_1108_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2235_ (.A1(_1120_),
    .A2(_0570_),
    .B(_0573_),
    .C(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2236_ (.A1(_0566_),
    .A2(_0577_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2237_ (.A1(_1187_),
    .A2(_1235_),
    .A3(_1245_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2238_ (.A1(_1205_),
    .A2(_1216_),
    .A3(_1217_),
    .A4(_1220_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2239_ (.A1(_1210_),
    .A2(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2240_ (.A1(_1202_),
    .A2(_1277_),
    .A3(_0579_),
    .A4(_0581_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2241_ (.I(\u1.ordering_timer[19] ),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2242_ (.A1(_0583_),
    .A2(_1058_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2243_ (.A1(_1062_),
    .A2(_1069_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2244_ (.A1(_1066_),
    .A2(_0585_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2245_ (.A1(_1051_),
    .A2(_1053_),
    .B(_1048_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2246_ (.A1(_1057_),
    .A2(_0584_),
    .A3(_0586_),
    .B1(_0587_),
    .B2(_1055_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2247_ (.A1(\u1.ordering_timer[27] ),
    .A2(_0506_),
    .B1(\u1.ordering_timer[26] ),
    .B2(_0504_),
    .C1(_1089_),
    .C2(_1092_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2248_ (.A1(_1084_),
    .A2(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2249_ (.I(_1080_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2250_ (.A1(_1077_),
    .A2(_0591_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2251_ (.A1(_1083_),
    .A2(_0592_),
    .B(_1074_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2252_ (.A1(_1095_),
    .A2(_0588_),
    .B(_0590_),
    .C(_0593_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2253_ (.A1(_1212_),
    .A2(_0578_),
    .A3(_0582_),
    .A4(_0594_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2254_ (.I(_0595_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2255_ (.I(_0596_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2256_ (.A1(_1139_),
    .A2(_0597_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2257_ (.A1(_0565_),
    .A2(_0598_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2258_ (.I(\u1.ordering_timer[1] ),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2259_ (.A1(_1403_),
    .A2(_0595_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2260_ (.I(_0600_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2261_ (.A1(_0565_),
    .A2(_0600_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2262_ (.I(_0602_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2263_ (.I(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2264_ (.A1(_1138_),
    .A2(_0599_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2265_ (.I(_0596_),
    .Z(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2266_ (.I(_0606_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2267_ (.I0(\u1.ordering_complete[1] ),
    .I1(_0605_),
    .S(_0607_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2268_ (.A1(_0599_),
    .A2(_0601_),
    .B1(_0604_),
    .B2(_0608_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2269_ (.I(_0609_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2270_ (.I(_0596_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2271_ (.I(_0610_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2272_ (.A1(_1138_),
    .A2(_0599_),
    .A3(\u1.ordering_timer[2] ),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2273_ (.A1(_1138_),
    .A2(_0599_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2274_ (.A1(_1136_),
    .A2(_0613_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2275_ (.A1(_0612_),
    .A2(_0614_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2276_ (.A1(\u1.ordering_complete[2] ),
    .A2(_0597_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2277_ (.A1(_0611_),
    .A2(_0615_),
    .B(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2278_ (.A1(\u1.ordering_timer[2] ),
    .A2(_0601_),
    .B1(_0604_),
    .B2(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2279_ (.I(_0618_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2280_ (.A1(\u1.ordering_timer[3] ),
    .A2(_0612_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2281_ (.A1(\u1.ordering_complete[3] ),
    .A2(_0597_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2282_ (.A1(_0611_),
    .A2(_0619_),
    .B(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2283_ (.A1(\u1.ordering_timer[3] ),
    .A2(_0601_),
    .B1(_0604_),
    .B2(_0621_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2284_ (.I(_0622_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2285_ (.I(\u1.ordering_timer[4] ),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2286_ (.I(_0600_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2287_ (.I(_0624_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2288_ (.I(_0625_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2289_ (.A1(\u1.ordering_timer[0] ),
    .A2(\u1.ordering_timer[1] ),
    .A3(\u1.ordering_timer[3] ),
    .A4(\u1.ordering_timer[2] ),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2290_ (.A1(_1122_),
    .A2(_0627_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2291_ (.I(_0595_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2292_ (.I(_0629_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2293_ (.A1(\u1.ordering_complete[4] ),
    .A2(_0630_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2294_ (.A1(_0611_),
    .A2(_0628_),
    .B(_0631_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2295_ (.A1(_0623_),
    .A2(_0626_),
    .B1(_0604_),
    .B2(_0632_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2296_ (.I(_0633_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2297_ (.I(_0602_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2298_ (.I(_0634_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2299_ (.A1(\u1.ordering_timer[5] ),
    .A2(_0623_),
    .A3(_0627_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2300_ (.A1(_0623_),
    .A2(_0627_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2301_ (.A1(_1121_),
    .A2(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2302_ (.A1(_0636_),
    .A2(_0638_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2303_ (.A1(\u1.ordering_complete[5] ),
    .A2(_0630_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2304_ (.A1(_0611_),
    .A2(_0639_),
    .B(_0640_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2305_ (.A1(\u1.ordering_timer[5] ),
    .A2(_0626_),
    .B1(_0635_),
    .B2(_0641_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2306_ (.I(_0642_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2307_ (.I(_0610_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2308_ (.A1(\u1.ordering_timer[6] ),
    .A2(_0636_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2309_ (.A1(\u1.ordering_complete[6] ),
    .A2(_0630_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2310_ (.A1(_0643_),
    .A2(_0644_),
    .B(_0645_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2311_ (.A1(\u1.ordering_timer[6] ),
    .A2(_0626_),
    .B1(_0635_),
    .B2(_0646_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2312_ (.I(_0647_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2313_ (.I(\u1.ordering_timer[7] ),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2314_ (.A1(\u1.ordering_timer[6] ),
    .A2(\u1.ordering_timer[5] ),
    .A3(_0623_),
    .A4(_0627_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2315_ (.A1(_1124_),
    .A2(_0649_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2316_ (.A1(\u1.ordering_complete[7] ),
    .A2(_0630_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2317_ (.A1(_0643_),
    .A2(_0650_),
    .B(_0651_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2318_ (.A1(_0648_),
    .A2(_0626_),
    .B1(_0635_),
    .B2(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2319_ (.I(_0653_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2320_ (.I(\u1.ordering_timer[8] ),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2321_ (.I(_0625_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2322_ (.A1(_0648_),
    .A2(_0649_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2323_ (.A1(_1111_),
    .A2(_0656_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2324_ (.I(_0629_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2325_ (.A1(_1112_),
    .A2(_0658_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2326_ (.A1(_0643_),
    .A2(_0657_),
    .B(_0659_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2327_ (.A1(_0654_),
    .A2(_0655_),
    .B1(_0635_),
    .B2(_0660_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2328_ (.I(_0661_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2329_ (.I(_0634_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2330_ (.A1(_0654_),
    .A2(_0656_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2331_ (.A1(_1109_),
    .A2(_0663_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2332_ (.A1(_0648_),
    .A2(\u1.ordering_timer[9] ),
    .A3(_0654_),
    .A4(_0649_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2333_ (.A1(_0664_),
    .A2(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2334_ (.A1(_1110_),
    .A2(_0658_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2335_ (.A1(_0643_),
    .A2(_0666_),
    .B(_0667_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2336_ (.A1(\u1.ordering_timer[9] ),
    .A2(_0655_),
    .B1(_0662_),
    .B2(_0668_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2337_ (.I(_0669_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2338_ (.I(_0610_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2339_ (.A1(\u1.ordering_timer[10] ),
    .A2(_0665_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2340_ (.A1(\u1.ordering_complete[10] ),
    .A2(_0658_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2341_ (.A1(_0670_),
    .A2(_0671_),
    .B(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2342_ (.A1(\u1.ordering_timer[10] ),
    .A2(_0655_),
    .B1(_0662_),
    .B2(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2343_ (.I(_0674_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2344_ (.I(\u1.ordering_timer[11] ),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2345_ (.I(_0675_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2346_ (.A1(_1116_),
    .A2(_0665_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2347_ (.A1(_0676_),
    .A2(_0677_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2348_ (.A1(\u1.ordering_complete[11] ),
    .A2(_0658_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2349_ (.A1(_0670_),
    .A2(_0678_),
    .B(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2350_ (.A1(_0675_),
    .A2(_0655_),
    .B1(_0662_),
    .B2(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2351_ (.I(_0681_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2352_ (.I(_0625_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2353_ (.A1(_0675_),
    .A2(_0677_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2354_ (.A1(_1103_),
    .A2(_0683_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2355_ (.A1(\u1.ordering_timer[12] ),
    .A2(_0675_),
    .A3(_0677_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2356_ (.A1(_0684_),
    .A2(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2357_ (.I(_0629_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2358_ (.A1(\u1.ordering_complete[12] ),
    .A2(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2359_ (.A1(_0670_),
    .A2(_0686_),
    .B(_0688_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2360_ (.A1(\u1.ordering_timer[12] ),
    .A2(_0682_),
    .B1(_0662_),
    .B2(_0689_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2361_ (.I(_0690_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2362_ (.I(_0634_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2363_ (.A1(\u1.ordering_timer[13] ),
    .A2(\u1.ordering_timer[12] ),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2364_ (.A1(_0676_),
    .A2(_1116_),
    .A3(_0665_),
    .A4(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2365_ (.I(_0693_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2366_ (.A1(_1101_),
    .A2(_0685_),
    .B(_0694_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2367_ (.I0(\u1.ordering_complete[13] ),
    .I1(_0695_),
    .S(_0607_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2368_ (.A1(\u1.ordering_timer[13] ),
    .A2(_0682_),
    .B1(_0691_),
    .B2(_0696_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2369_ (.I(_0697_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2370_ (.I(\u1.ordering_timer[14] ),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2371_ (.A1(_1100_),
    .A2(_0694_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2372_ (.A1(\u1.ordering_complete[14] ),
    .A2(_0687_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2373_ (.A1(_0670_),
    .A2(_0699_),
    .B(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2374_ (.A1(_0698_),
    .A2(_0682_),
    .B1(_0691_),
    .B2(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2375_ (.I(_0702_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2376_ (.I(_1096_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2377_ (.A1(_0698_),
    .A2(_0694_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2378_ (.A1(_0703_),
    .A2(_0704_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2379_ (.I0(\u1.ordering_complete[15] ),
    .I1(_0705_),
    .S(_0607_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2380_ (.A1(_0703_),
    .A2(_0682_),
    .B1(_0691_),
    .B2(_0706_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2381_ (.I(_0707_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2382_ (.I(_1059_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2383_ (.I(_0624_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2384_ (.I(_0709_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2385_ (.I(_0606_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2386_ (.A1(_0703_),
    .A2(_0698_),
    .A3(_0694_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2387_ (.A1(_1059_),
    .A2(_0712_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2388_ (.I(_0606_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2389_ (.A1(\u1.ordering_complete[16] ),
    .A2(_0714_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2390_ (.I(_0624_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2391_ (.A1(_0711_),
    .A2(_0713_),
    .B(_0715_),
    .C(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2392_ (.A1(_0329_),
    .A2(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2393_ (.A1(_0708_),
    .A2(_0710_),
    .B(_0718_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2394_ (.I(_0625_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2395_ (.I(_0610_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2396_ (.A1(_0708_),
    .A2(_0712_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2397_ (.A1(_1068_),
    .A2(_1059_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2398_ (.A1(_1096_),
    .A2(\u1.ordering_timer[14] ),
    .A3(_0693_),
    .A4(_0722_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2399_ (.I(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2400_ (.I(_0596_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2401_ (.A1(_1068_),
    .A2(_0721_),
    .B(_0724_),
    .C(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2402_ (.A1(_1061_),
    .A2(_0720_),
    .B(_0726_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2403_ (.A1(_1068_),
    .A2(_0719_),
    .B1(_0691_),
    .B2(_0727_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2404_ (.I(_0728_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2405_ (.I(_1065_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2406_ (.A1(_0729_),
    .A2(_0723_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2407_ (.A1(\u1.ordering_complete[18] ),
    .A2(_0725_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2408_ (.A1(_0711_),
    .A2(_0730_),
    .B(_0731_),
    .C(_0716_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2409_ (.A1(_0329_),
    .A2(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2410_ (.A1(_0729_),
    .A2(_0710_),
    .B(_0733_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2411_ (.I(_0634_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2412_ (.I(_0606_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2413_ (.A1(\u1.ordering_timer[18] ),
    .A2(_0723_),
    .B(_0583_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2414_ (.A1(_1064_),
    .A2(_0729_),
    .A3(_0724_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2415_ (.A1(_0736_),
    .A2(_0737_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2416_ (.A1(\u1.ordering_complete[19] ),
    .A2(_0687_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2417_ (.A1(_0735_),
    .A2(_0738_),
    .B(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2418_ (.A1(_0583_),
    .A2(_0719_),
    .B1(_0734_),
    .B2(_0740_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2419_ (.I(_0741_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2420_ (.A1(_1050_),
    .A2(_0737_),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2421_ (.A1(\u1.ordering_complete[20] ),
    .A2(_0687_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2422_ (.A1(_0735_),
    .A2(_0742_),
    .B(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2423_ (.A1(\u1.ordering_timer[20] ),
    .A2(_0719_),
    .B1(_0734_),
    .B2(_0744_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2424_ (.I(_0745_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2425_ (.A1(\u1.ordering_timer[20] ),
    .A2(_0737_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2426_ (.A1(\u1.ordering_timer[21] ),
    .A2(\u1.ordering_timer[20] ),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2427_ (.I(_0747_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2428_ (.A1(_0583_),
    .A2(\u1.ordering_timer[18] ),
    .A3(_0723_),
    .A4(_0748_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2429_ (.I(_0749_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2430_ (.A1(_1049_),
    .A2(_0746_),
    .B(_0750_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2431_ (.I0(\u1.ordering_complete[21] ),
    .I1(_0751_),
    .S(_0714_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2432_ (.A1(\u1.ordering_timer[21] ),
    .A2(_0719_),
    .B1(_0734_),
    .B2(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2433_ (.I(_0753_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2434_ (.I(\u1.ordering_timer[22] ),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2435_ (.I(_0624_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2436_ (.A1(_1047_),
    .A2(_0750_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2437_ (.I(_0629_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2438_ (.A1(\u1.ordering_complete[22] ),
    .A2(_0757_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2439_ (.A1(_0735_),
    .A2(_0756_),
    .B(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2440_ (.A1(_0754_),
    .A2(_0755_),
    .B1(_0734_),
    .B2(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2441_ (.I(_0760_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2442_ (.I(\u1.ordering_timer[23] ),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2443_ (.I(_0602_),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2444_ (.A1(_0754_),
    .A2(_0750_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2445_ (.A1(_1046_),
    .A2(_0763_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2446_ (.A1(_0761_),
    .A2(_0754_),
    .A3(_0750_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2447_ (.A1(_0757_),
    .A2(_0764_),
    .A3(_0765_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2448_ (.A1(_1054_),
    .A2(_0720_),
    .B(_0766_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2449_ (.A1(_0761_),
    .A2(_0755_),
    .B1(_0762_),
    .B2(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2450_ (.I(_0768_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2451_ (.I(_1085_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2452_ (.A1(_0769_),
    .A2(_0765_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2453_ (.A1(\u1.ordering_complete[24] ),
    .A2(_0757_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2454_ (.A1(_0735_),
    .A2(_0770_),
    .B(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2455_ (.A1(_0769_),
    .A2(_0755_),
    .B1(_0762_),
    .B2(_0772_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2456_ (.I(_0773_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2457_ (.I(\u1.ordering_timer[25] ),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2458_ (.A1(_0648_),
    .A2(\u1.ordering_timer[9] ),
    .A3(_0654_),
    .A4(_0649_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2459_ (.A1(_0676_),
    .A2(_1116_),
    .A3(_0775_),
    .A4(_0692_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2460_ (.A1(_0703_),
    .A2(_0698_),
    .A3(_0776_),
    .A4(_0722_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2461_ (.A1(_1064_),
    .A2(_0729_),
    .A3(_0777_),
    .A4(_0747_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2462_ (.A1(_1085_),
    .A2(_0761_),
    .A3(_0754_),
    .A4(_0778_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2463_ (.A1(_0774_),
    .A2(_0779_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2464_ (.I0(\u1.ordering_complete[25] ),
    .I1(_0780_),
    .S(_0714_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2465_ (.A1(_0774_),
    .A2(_0755_),
    .B1(_0762_),
    .B2(_0781_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2466_ (.I(_0782_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2467_ (.I(\u1.ordering_timer[26] ),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2468_ (.A1(_0774_),
    .A2(_0761_),
    .A3(\u1.ordering_timer[22] ),
    .A4(_0749_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2469_ (.A1(_0769_),
    .A2(_0784_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2470_ (.A1(_1087_),
    .A2(_0785_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2471_ (.A1(\u1.ordering_complete[26] ),
    .A2(_0757_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2472_ (.A1(_0711_),
    .A2(_0786_),
    .B(_0787_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2473_ (.A1(_0783_),
    .A2(_0716_),
    .B1(_0762_),
    .B2(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2474_ (.I(_0789_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2475_ (.A1(_0783_),
    .A2(_0774_),
    .A3(_0779_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2476_ (.A1(\u1.ordering_timer[27] ),
    .A2(_0783_),
    .A3(_1085_),
    .A4(_0784_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2477_ (.I(_0725_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2478_ (.A1(_1093_),
    .A2(_0790_),
    .B(_0791_),
    .C(_0792_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2479_ (.A1(_0506_),
    .A2(_0711_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2480_ (.A1(_0793_),
    .A2(_0794_),
    .B(_0603_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2481_ (.A1(_1093_),
    .A2(_0710_),
    .B(_0795_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2482_ (.I(_1071_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2483_ (.A1(_0796_),
    .A2(_0791_),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2484_ (.A1(_0597_),
    .A2(_0797_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2485_ (.A1(\u1.ordering_complete[28] ),
    .A2(_0720_),
    .B(_0603_),
    .C(_0798_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2486_ (.A1(_0796_),
    .A2(_0710_),
    .B(_0799_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2487_ (.A1(\u1.ordering_timer[28] ),
    .A2(_0791_),
    .B(\u1.ordering_timer[29] ),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2488_ (.A1(_1076_),
    .A2(_0796_),
    .A3(_1093_),
    .A4(_0790_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2489_ (.A1(_0800_),
    .A2(_0801_),
    .B(_0607_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2490_ (.A1(\u1.ordering_complete[29] ),
    .A2(_0720_),
    .B(_0709_),
    .C(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2491_ (.A1(_1076_),
    .A2(_0709_),
    .B1(_0803_),
    .B2(_0565_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2492_ (.A1(\u1.ordering_complete[30] ),
    .A2(_0792_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2493_ (.A1(_1082_),
    .A2(\u1.ordering_timer[29] ),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2494_ (.A1(\u1.ordering_timer[28] ),
    .A2(_0791_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2495_ (.A1(_1082_),
    .A2(_0801_),
    .B1(_0805_),
    .B2(_0806_),
    .C(_0725_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2496_ (.A1(_0804_),
    .A2(_0807_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2497_ (.A1(_1082_),
    .A2(_0716_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2498_ (.A1(_0565_),
    .A2(_0601_),
    .A3(_0808_),
    .B(_0809_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2499_ (.I(\u1.ordering_timer[31] ),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2500_ (.A1(\u1.ordering_timer[27] ),
    .A2(_0783_),
    .A3(_0769_),
    .A4(_0784_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2501_ (.A1(_0796_),
    .A2(_0811_),
    .A3(_0805_),
    .B(_0810_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2502_ (.I0(\u1.ordering_complete[31] ),
    .I1(_0812_),
    .S(_0714_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2503_ (.A1(_0603_),
    .A2(_0813_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2504_ (.A1(_0810_),
    .A2(_0709_),
    .B(_0814_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2505_ (.I(_1041_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2506_ (.A1(_0815_),
    .A2(\u0.latch_cmd ),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2507_ (.I(_0816_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2508_ (.I(_0817_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2509_ (.A1(_1042_),
    .A2(\u0.latch_cmd ),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2510_ (.I(_0819_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2511_ (.I(_0820_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2512_ (.A1(_0513_),
    .A2(_0818_),
    .B1(_0821_),
    .B2(\spi_data_crossing[0].data_sync ),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2513_ (.I(_0822_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2514_ (.A1(_0517_),
    .A2(_0818_),
    .B1(_0821_),
    .B2(\spi_data_crossing[1].data_sync ),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2515_ (.I(_0823_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2516_ (.A1(_0459_),
    .A2(_0818_),
    .B1(_0821_),
    .B2(\spi_data_crossing[2].data_sync ),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2517_ (.I(_0824_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2518_ (.A1(_0462_),
    .A2(_0818_),
    .B1(_0821_),
    .B2(\spi_data_crossing[3].data_sync ),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2519_ (.I(_0825_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2520_ (.I(_0817_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2521_ (.I(_0820_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2522_ (.A1(_0464_),
    .A2(_0826_),
    .B1(_0827_),
    .B2(\spi_data_crossing[4].data_sync ),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2523_ (.I(_0828_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2524_ (.A1(_0466_),
    .A2(_0826_),
    .B1(_0827_),
    .B2(\spi_data_crossing[5].data_sync ),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2525_ (.I(_0829_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2526_ (.A1(_0469_),
    .A2(_0826_),
    .B1(_0827_),
    .B2(\spi_data_crossing[6].data_sync ),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2527_ (.I(_0830_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2528_ (.A1(_0472_),
    .A2(_0826_),
    .B1(_0827_),
    .B2(\spi_data_crossing[7].data_sync ),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2529_ (.I(_0831_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2530_ (.I(_0817_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2531_ (.I(_0820_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2532_ (.A1(_0474_),
    .A2(_0832_),
    .B1(_0833_),
    .B2(\spi_data_crossing[8].data_sync ),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2533_ (.I(_0834_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2534_ (.A1(_0476_),
    .A2(_0832_),
    .B1(_0833_),
    .B2(\spi_data_crossing[9].data_sync ),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2535_ (.I(_0835_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2536_ (.A1(_0379_),
    .A2(_0832_),
    .B1(_0833_),
    .B2(\spi_data_crossing[10].data_sync ),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2537_ (.I(_0836_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2538_ (.A1(_0381_),
    .A2(_0832_),
    .B1(_0833_),
    .B2(\spi_data_crossing[11].data_sync ),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2539_ (.I(_0837_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2540_ (.I(_0817_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2541_ (.I(_0820_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2542_ (.A1(_0442_),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\spi_data_crossing[12].data_sync ),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2543_ (.I(_0840_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2544_ (.A1(_0385_),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\spi_data_crossing[13].data_sync ),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2545_ (.I(_0841_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2546_ (.A1(_0387_),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\spi_data_crossing[14].data_sync ),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2547_ (.I(_0842_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2548_ (.A1(_0389_),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\spi_data_crossing[15].data_sync ),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2549_ (.I(_0843_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2550_ (.I(_0816_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2551_ (.I(_0844_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2552_ (.I(_0819_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2553_ (.I(_0846_),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2554_ (.A1(_0447_),
    .A2(_0845_),
    .B1(_0847_),
    .B2(\spi_data_crossing[16].data_sync ),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2555_ (.I(_0848_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2556_ (.A1(_0348_),
    .A2(_0845_),
    .B1(_0847_),
    .B2(\spi_data_crossing[17].data_sync ),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2557_ (.I(_0849_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2558_ (.A1(\u0.cmd[18] ),
    .A2(_0845_),
    .B1(_0847_),
    .B2(\spi_data_crossing[18].data_sync ),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2559_ (.I(_0850_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2560_ (.A1(\u0.cmd[19] ),
    .A2(_0845_),
    .B1(_0847_),
    .B2(\spi_data_crossing[19].data_sync ),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2561_ (.I(_0851_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2562_ (.I(_0844_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2563_ (.I(_0846_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2564_ (.A1(\u0.cmd[20] ),
    .A2(_0852_),
    .B1(_0853_),
    .B2(\spi_data_crossing[20].data_sync ),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2565_ (.I(_0854_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2566_ (.A1(\u0.cmd[21] ),
    .A2(_0852_),
    .B1(_0853_),
    .B2(\spi_data_crossing[21].data_sync ),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2567_ (.I(_0855_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2568_ (.A1(\u0.cmd[22] ),
    .A2(_0852_),
    .B1(_0853_),
    .B2(\spi_data_crossing[22].data_sync ),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2569_ (.I(_0856_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2570_ (.A1(\u0.cmd[23] ),
    .A2(_0852_),
    .B1(_0853_),
    .B2(\spi_data_crossing[23].data_sync ),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2571_ (.I(_0857_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2572_ (.I(_0844_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2573_ (.I(_0846_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2574_ (.A1(\u0.cmd[24] ),
    .A2(_0858_),
    .B1(_0859_),
    .B2(\spi_data_crossing[24].data_sync ),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2575_ (.I(_0860_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2576_ (.A1(\u0.cmd[25] ),
    .A2(_0858_),
    .B1(_0859_),
    .B2(\spi_data_crossing[25].data_sync ),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2577_ (.I(_0861_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2578_ (.A1(_0299_),
    .A2(_0858_),
    .B1(_0859_),
    .B2(\spi_data_crossing[26].data_sync ),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2579_ (.I(_0862_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2580_ (.A1(_1160_),
    .A2(_0858_),
    .B1(_0859_),
    .B2(\spi_data_crossing[27].data_sync ),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2581_ (.I(_0863_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2582_ (.I(_0844_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2583_ (.I(_0846_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2584_ (.A1(\u0.cmd[28] ),
    .A2(_0864_),
    .B1(_0865_),
    .B2(\spi_data_crossing[28].data_sync ),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2585_ (.I(_0866_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2586_ (.A1(_1153_),
    .A2(_0864_),
    .B1(_0865_),
    .B2(\spi_data_crossing[29].data_sync ),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2587_ (.I(_0867_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2588_ (.A1(\u0.cmd[30] ),
    .A2(_0864_),
    .B1(_0865_),
    .B2(\spi_data_crossing[30].data_sync ),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2589_ (.I(_0868_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2590_ (.A1(_1040_),
    .A2(_0864_),
    .B1(_0865_),
    .B2(\spi_data_crossing[31].data_sync ),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2591_ (.I(_0869_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2592_ (.A1(\u1.col_sel[0] ),
    .A2(_0321_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2593_ (.A1(_0312_),
    .A2(_0324_),
    .A3(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2594_ (.A1(_0322_),
    .A2(_0326_),
    .A3(_0871_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2595_ (.A1(_0313_),
    .A2(\u1.col_limit[3] ),
    .B1(_0316_),
    .B2(\u1.col_limit[2] ),
    .C(_0315_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2596_ (.A1(_0320_),
    .A2(_0872_),
    .A3(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2597_ (.A1(_0309_),
    .A2(_0874_),
    .B(_1212_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2598_ (.I(\u1.row_sel[4] ),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2599_ (.I(\u1.row_sel[3] ),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2600_ (.I(\u1.row_sel[1] ),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2601_ (.I(\u1.row_sel[0] ),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2602_ (.A1(\u1.row_limit[1] ),
    .A2(_0878_),
    .B(\u1.row_limit[0] ),
    .C(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2603_ (.I(\u1.row_sel[2] ),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2604_ (.A1(\u1.row_limit[2] ),
    .A2(_0881_),
    .B1(\u1.row_limit[1] ),
    .B2(_0878_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2605_ (.A1(\u1.row_limit[3] ),
    .A2(_0877_),
    .B1(\u1.row_limit[2] ),
    .B2(_0881_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2606_ (.A1(_0880_),
    .A2(_0882_),
    .B(_0883_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2607_ (.A1(\u1.row_limit[4] ),
    .A2(_0876_),
    .B1(\u1.row_limit[3] ),
    .B2(_0877_),
    .C(_0884_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2608_ (.A1(_0524_),
    .A2(\u1.row_sel[5] ),
    .B1(_0521_),
    .B2(\u1.row_sel[4] ),
    .C(_0885_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2609_ (.A1(\u1.row_sel[6] ),
    .A2(_0526_),
    .B1(_0524_),
    .B2(\u1.row_sel[5] ),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2610_ (.A1(\u1.row_sel[6] ),
    .A2(_0526_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2611_ (.A1(_0886_),
    .A2(_0887_),
    .B(_0888_),
    .C(_0329_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2612_ (.A1(_0875_),
    .A2(_0889_),
    .Z(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2613_ (.I(_0890_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2614_ (.A1(\u1.row_sel[0] ),
    .A2(_0875_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2615_ (.A1(\u1.row_sel[0] ),
    .A2(_0875_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2616_ (.A1(_0891_),
    .A2(_0892_),
    .A3(_0893_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2617_ (.A1(_0878_),
    .A2(_0892_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2618_ (.A1(_0891_),
    .A2(_0894_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2619_ (.A1(\u1.row_sel[2] ),
    .A2(\u1.row_sel[1] ),
    .A3(_0892_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2620_ (.A1(\u1.row_sel[1] ),
    .A2(_0892_),
    .B(\u1.row_sel[2] ),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2621_ (.A1(_0890_),
    .A2(_0895_),
    .A3(_0896_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2622_ (.A1(\u1.row_sel[3] ),
    .A2(_0895_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2623_ (.A1(\u1.row_sel[3] ),
    .A2(_0895_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2624_ (.A1(_0890_),
    .A2(_0897_),
    .A3(_0898_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2625_ (.A1(\u1.row_sel[4] ),
    .A2(_0897_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2626_ (.A1(\u1.row_sel[4] ),
    .A2(_0897_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2627_ (.A1(_0890_),
    .A2(_0899_),
    .A3(_0900_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2628_ (.I(\u1.row_sel[5] ),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2629_ (.A1(_0901_),
    .A2(_0900_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2630_ (.A1(_0891_),
    .A2(_0902_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2631_ (.A1(\u1.row_sel[5] ),
    .A2(_0900_),
    .B(\u1.row_sel[6] ),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2632_ (.A1(_0891_),
    .A2(_0903_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2633_ (.A1(\latch_data_sync[0] ),
    .A2(latch_data),
    .A3(\latch_data_sync[1] ),
    .A4(_1042_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2634_ (.I(_0904_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2635_ (.A1(_1156_),
    .A2(_0815_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2636_ (.I(net20),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2637_ (.A1(_0905_),
    .A2(net38),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2638_ (.A1(\u1.ccr1[11] ),
    .A2(_1269_),
    .B1(\u1.ccr1[10] ),
    .B2(_1268_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2639_ (.A1(_0906_),
    .A2(_1270_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2640_ (.A1(_1274_),
    .A2(_1251_),
    .A3(_1275_),
    .B(_0907_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2641_ (.A1(_1252_),
    .A2(_1303_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2642_ (.A1(_1255_),
    .A2(_0909_),
    .B1(_1260_),
    .B2(_1264_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2643_ (.A1(\u1.ccr1[7] ),
    .A2(_1193_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2644_ (.A1(_1200_),
    .A2(_1188_),
    .B1(_1196_),
    .B2(_1190_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2645_ (.A1(_0912_),
    .A2(_1198_),
    .B(_1201_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2646_ (.A1(_1210_),
    .A2(_1218_),
    .B(_1205_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2647_ (.A1(_1216_),
    .A2(_0914_),
    .B(_1219_),
    .C(_1202_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2648_ (.A1(_0911_),
    .A2(_0913_),
    .B(_0915_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2649_ (.A1(_1277_),
    .A2(_0916_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2650_ (.A1(_1266_),
    .A2(_0908_),
    .B(_0910_),
    .C(_0917_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2651_ (.A1(_1227_),
    .A2(_1231_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2652_ (.A1(_0429_),
    .A2(_1318_),
    .B(_1321_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2653_ (.A1(_1241_),
    .A2(_1238_),
    .A3(_1242_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2654_ (.A1(_0429_),
    .A2(\u1.timer[19] ),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2655_ (.A1(\u1.ccr1[18] ),
    .A2(_0920_),
    .B(_0921_),
    .C(_0922_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2656_ (.A1(\u1.ccr1[23] ),
    .A2(_1228_),
    .B(_1227_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2657_ (.A1(_0919_),
    .A2(_1234_),
    .B1(_1235_),
    .B2(_0923_),
    .C(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2658_ (.A1(_1246_),
    .A2(_0918_),
    .B(_0925_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2659_ (.A1(_1187_),
    .A2(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2660_ (.A1(\u1.ccr1[25] ),
    .A2(_1164_),
    .B1(\u1.ccr1[24] ),
    .B2(_1166_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2661_ (.A1(_0928_),
    .A2(_1181_),
    .A3(_1183_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2662_ (.A1(\u1.ccr1[28] ),
    .A2(_1173_),
    .B1(\u1.ccr1[27] ),
    .B2(_1349_),
    .C1(_1179_),
    .C2(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2663_ (.A1(_1169_),
    .A2(_1172_),
    .B1(_1175_),
    .B2(_0930_),
    .C(_1185_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2664_ (.A1(_1402_),
    .A2(_0927_),
    .A3(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2665_ (.A1(_1279_),
    .A2(_0932_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2666_ (.I(_0933_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2667_ (.I(_0934_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2668_ (.A1(_1206_),
    .A2(_0935_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2669_ (.A1(_1364_),
    .A2(_1208_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2670_ (.A1(_0935_),
    .A2(_0936_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2671_ (.I(_0933_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2672_ (.A1(_1364_),
    .A2(_1363_),
    .A3(_1204_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2673_ (.A1(_1206_),
    .A2(_1208_),
    .B(_1203_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2674_ (.A1(_0937_),
    .A2(_0938_),
    .A3(_0939_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2675_ (.A1(_1214_),
    .A2(_0938_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2676_ (.A1(\u1.timer[0] ),
    .A2(\u1.timer[1] ),
    .A3(\u1.timer[3] ),
    .A4(\u1.timer[2] ),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2677_ (.A1(_0937_),
    .A2(_0940_),
    .A3(_0941_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2678_ (.A1(_1287_),
    .A2(_0941_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2679_ (.A1(_1287_),
    .A2(_0941_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2680_ (.A1(_0937_),
    .A2(_0942_),
    .A3(_0943_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2681_ (.A1(_1191_),
    .A2(_0942_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2682_ (.A1(_0935_),
    .A2(_0944_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2683_ (.I(_0933_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2684_ (.I(_0945_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2685_ (.A1(\u1.timer[6] ),
    .A2(\u1.timer[5] ),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2686_ (.A1(_0942_),
    .A2(_0947_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2687_ (.A1(_1283_),
    .A2(_0942_),
    .B(_1280_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2688_ (.A1(_0946_),
    .A2(_0948_),
    .A3(_0949_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2689_ (.A1(\u1.timer[7] ),
    .A2(\u1.timer[4] ),
    .A3(_0941_),
    .A4(_0947_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2690_ (.I(_0950_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2691_ (.A1(_1289_),
    .A2(_0948_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2692_ (.A1(_0946_),
    .A2(_0951_),
    .A3(_0952_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2693_ (.A1(_1250_),
    .A2(_0951_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2694_ (.A1(_1250_),
    .A2(_0951_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2695_ (.A1(_0946_),
    .A2(_0953_),
    .A3(_0954_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2696_ (.A1(_1293_),
    .A2(_1267_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2697_ (.A1(_0951_),
    .A2(_0955_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2698_ (.A1(_1248_),
    .A2(_0954_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2699_ (.A1(_0946_),
    .A2(_0956_),
    .A3(_0957_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2700_ (.I(_0945_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2701_ (.A1(_1295_),
    .A2(_0956_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2702_ (.A1(_1295_),
    .A2(_0956_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2703_ (.A1(_0958_),
    .A2(_0959_),
    .A3(_0960_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2704_ (.A1(_1272_),
    .A2(\u1.timer[10] ),
    .A3(_0950_),
    .A4(_0955_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2705_ (.A1(_1272_),
    .A2(_0959_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2706_ (.A1(_0958_),
    .A2(_0961_),
    .A3(_0962_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2707_ (.A1(_1311_),
    .A2(_0961_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2708_ (.A1(_1311_),
    .A2(_0961_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2709_ (.A1(_0958_),
    .A2(_0963_),
    .A3(_0964_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2710_ (.A1(_1258_),
    .A2(_0963_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2711_ (.A1(_0935_),
    .A2(_0965_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2712_ (.A1(_1254_),
    .A2(_1300_),
    .A3(_1262_),
    .A4(_0961_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2713_ (.A1(_1300_),
    .A2(_0963_),
    .B(_1254_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2714_ (.A1(_0958_),
    .A2(_0966_),
    .A3(_0967_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2715_ (.I(_0945_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2716_ (.A1(_1303_),
    .A2(_0966_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2717_ (.A1(_1303_),
    .A2(_0966_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2718_ (.I(_0970_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2719_ (.A1(_0968_),
    .A2(_0969_),
    .A3(_0971_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2720_ (.A1(_0283_),
    .A2(_0971_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2721_ (.A1(_1279_),
    .A2(_0932_),
    .B1(_0971_),
    .B2(_0283_),
    .C(_0972_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2722_ (.A1(_0283_),
    .A2(_0971_),
    .B(_0282_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2723_ (.A1(_0282_),
    .A2(\u1.timer[16] ),
    .A3(_0970_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2724_ (.A1(_0968_),
    .A2(_0973_),
    .A3(_0974_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2725_ (.A1(_1322_),
    .A2(_0974_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2726_ (.A1(_1321_),
    .A2(_0282_),
    .A3(\u1.timer[16] ),
    .A4(_0970_),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2727_ (.A1(_0968_),
    .A2(_0975_),
    .A3(_0976_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2728_ (.A1(_0281_),
    .A2(_0976_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2729_ (.A1(_0281_),
    .A2(_1322_),
    .A3(_0974_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2730_ (.A1(_0968_),
    .A2(_0977_),
    .A3(_0978_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2731_ (.A1(_1224_),
    .A2(_0978_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2732_ (.A1(_0937_),
    .A2(_0979_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2733_ (.A1(\u1.timer[20] ),
    .A2(_0978_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2734_ (.A1(\u1.timer[21] ),
    .A2(\u1.timer[20] ),
    .A3(_0281_),
    .A4(_0976_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2735_ (.I(_0933_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2736_ (.A1(_1233_),
    .A2(_0980_),
    .B(_0981_),
    .C(_0982_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2737_ (.I(_0945_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2738_ (.A1(_0286_),
    .A2(_0981_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2739_ (.A1(_0286_),
    .A2(_0981_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2740_ (.A1(_0983_),
    .A2(_0984_),
    .A3(_0985_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2741_ (.A1(_0285_),
    .A2(_0985_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2742_ (.A1(_0285_),
    .A2(_0985_),
    .B(_0986_),
    .C(_0982_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2743_ (.A1(_0285_),
    .A2(_0985_),
    .B(\u1.timer[24] ),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2744_ (.A1(\u1.timer[24] ),
    .A2(_1327_),
    .A3(_0286_),
    .A4(_0981_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2745_ (.A1(_0983_),
    .A2(_0987_),
    .A3(_0988_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2746_ (.A1(_1411_),
    .A2(_0988_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2747_ (.A1(_1411_),
    .A2(_0988_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2748_ (.A1(_0983_),
    .A2(_0989_),
    .A3(_0990_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2749_ (.A1(_1410_),
    .A2(_0990_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2750_ (.A1(_1410_),
    .A2(_0990_),
    .B(_0991_),
    .C(_0982_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2751_ (.A1(_1410_),
    .A2(_0990_),
    .B(_1394_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2752_ (.A1(_1394_),
    .A2(_1345_),
    .A3(_1411_),
    .A4(_0988_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2753_ (.A1(_0983_),
    .A2(_0992_),
    .A3(_0993_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2754_ (.A1(_1413_),
    .A2(_0993_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2755_ (.A1(_1413_),
    .A2(_0993_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2756_ (.A1(_0982_),
    .A2(_0994_),
    .A3(_0995_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2757_ (.I(\u1.timer[29] ),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2758_ (.A1(_0996_),
    .A2(_0995_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2759_ (.A1(_0996_),
    .A2(_0995_),
    .B(_0997_),
    .C(_0934_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2760_ (.A1(_0996_),
    .A2(_0995_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2761_ (.A1(\u1.timer[30] ),
    .A2(_0996_),
    .A3(_1413_),
    .A4(_0993_),
    .Z(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2762_ (.A1(_1167_),
    .A2(_0998_),
    .B(_0999_),
    .C(_0934_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2763_ (.A1(_1351_),
    .A2(_0999_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2764_ (.A1(_1351_),
    .A2(_0999_),
    .B(_1000_),
    .C(_0934_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2765_ (.I(net12),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2766_ (.A1(_1001_),
    .A2(net30),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2767_ (.I(net11),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2768_ (.A1(_1002_),
    .A2(net29),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2769_ (.I(net10),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2770_ (.A1(_1003_),
    .A2(net28),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2771_ (.I(net9),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2772_ (.A1(_1004_),
    .A2(net27),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2773_ (.I(net8),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2774_ (.A1(_1005_),
    .A2(net26),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2775_ (.I(net7),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2776_ (.A1(_1006_),
    .A2(net25),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2777_ (.I(net6),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2778_ (.A1(_1007_),
    .A2(net24),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2779_ (.I(net5),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2780_ (.A1(_1008_),
    .A2(net23),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2781_ (.I(net21),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2782_ (.A1(_1009_),
    .A2(net39),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2783_ (.I(\u1.ccr0[0] ),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2784_ (.A1(_0447_),
    .A2(_0347_),
    .A3(_0351_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2785_ (.I(_1011_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2786_ (.I(_1012_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2787_ (.I(_1013_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2788_ (.I(_1012_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2789_ (.A1(_0345_),
    .A2(_1015_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2790_ (.A1(_1010_),
    .A2(_1014_),
    .B(_1016_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2791_ (.I(_1012_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2792_ (.I0(\u1.ccr0[1] ),
    .I1(_0356_),
    .S(_1017_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2793_ (.I(_1018_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2794_ (.I0(\u1.ccr0[2] ),
    .I1(_0360_),
    .S(_1017_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2795_ (.I(_1019_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2796_ (.I0(\u1.ccr0[3] ),
    .I1(_0363_),
    .S(_1013_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2797_ (.I(_1020_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2798_ (.I(_1011_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2799_ (.A1(_0404_),
    .A2(_1021_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2800_ (.A1(_1286_),
    .A2(_1014_),
    .B(_1022_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2801_ (.A1(_0406_),
    .A2(_1021_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2802_ (.A1(_1282_),
    .A2(_1014_),
    .B(_1023_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2803_ (.A1(_0468_),
    .A2(_1021_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2804_ (.A1(_1281_),
    .A2(_1014_),
    .B(_1024_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2805_ (.I(_1012_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2806_ (.A1(_0372_),
    .A2(_1021_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2807_ (.A1(_1290_),
    .A2(_1025_),
    .B(_1026_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2808_ (.I0(\u1.ccr0[8] ),
    .I1(_0374_),
    .S(_1013_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2809_ (.I(_1027_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2810_ (.I0(\u1.ccr0[9] ),
    .I1(_0376_),
    .S(_1013_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2811_ (.I(_1028_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2812_ (.I(_1011_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2813_ (.A1(\u0.cmd[10] ),
    .A2(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2814_ (.A1(_1296_),
    .A2(_1025_),
    .B(_1030_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2815_ (.I(\u1.ccr0[11] ),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2816_ (.A1(\u0.cmd[11] ),
    .A2(_1029_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2817_ (.A1(_1031_),
    .A2(_1025_),
    .B(_1032_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2818_ (.A1(\u0.cmd[12] ),
    .A2(_1029_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2819_ (.A1(_1310_),
    .A2(_1025_),
    .B(_1033_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2820_ (.A1(\u0.cmd[13] ),
    .A2(_1029_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2821_ (.A1(_1301_),
    .A2(_1015_),
    .B(_1034_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2822_ (.A1(\u0.cmd[14] ),
    .A2(_1017_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2823_ (.A1(_1305_),
    .A2(_1015_),
    .B(_1035_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2824_ (.A1(\u0.cmd[15] ),
    .A2(_1017_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2825_ (.A1(_1304_),
    .A2(_1015_),
    .B(_1036_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2826_ (.A1(net4),
    .A2(net22),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2827_ (.I(_1037_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2828_ (.A1(net13),
    .A2(net31),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2829_ (.I(_1038_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2830_ (.A1(net14),
    .A2(net32),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2831_ (.I(_1039_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2832_ (.D(\u1.row_sel[0] ),
    .CLK(clknet_leaf_13_clock),
    .Q(net204));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2833_ (.D(\u1.row_sel[1] ),
    .CLK(clknet_leaf_13_clock),
    .Q(net205));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2834_ (.D(\u1.row_sel[2] ),
    .CLK(clknet_leaf_13_clock),
    .Q(net206));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2835_ (.D(\u1.row_sel[3] ),
    .CLK(clknet_leaf_13_clock),
    .Q(net207));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2836_ (.D(\u1.row_sel[4] ),
    .CLK(clknet_leaf_13_clock),
    .Q(net208));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2837_ (.D(\u1.row_sel[5] ),
    .CLK(clknet_leaf_13_clock),
    .Q(net209));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2838_ (.D(\u1.col_sel[0] ),
    .CLK(clknet_leaf_18_clock),
    .Q(net83));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2839_ (.D(\u1.col_sel[1] ),
    .CLK(clknet_leaf_18_clock),
    .Q(net84));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2840_ (.D(\u1.col_sel[2] ),
    .CLK(clknet_leaf_18_clock),
    .Q(net85));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2841_ (.D(\u1.col_sel[3] ),
    .CLK(clknet_leaf_19_clock),
    .Q(net86));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2842_ (.D(\u1.col_sel[4] ),
    .CLK(clknet_leaf_19_clock),
    .Q(net87));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2843_ (.D(\u1.col_sel[5] ),
    .CLK(clknet_leaf_19_clock),
    .Q(net88));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2844_ (.D(\u0.cmd[0] ),
    .CLK(clknet_leaf_17_clock),
    .Q(net95));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2845_ (.D(\u0.cmd[1] ),
    .CLK(clknet_leaf_18_clock),
    .Q(net102));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2846_ (.D(\u0.cmd[2] ),
    .CLK(clknet_leaf_17_clock),
    .Q(net103));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2847_ (.D(\u0.cmd[3] ),
    .CLK(clknet_leaf_19_clock),
    .Q(net104));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2848_ (.D(\u0.cmd[4] ),
    .CLK(clknet_leaf_23_clock),
    .Q(net105));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2849_ (.D(\u0.cmd[5] ),
    .CLK(clknet_leaf_20_clock),
    .Q(net106));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2850_ (.D(\u0.cmd[6] ),
    .CLK(clknet_leaf_20_clock),
    .Q(net107));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2851_ (.D(\u0.cmd[7] ),
    .CLK(clknet_leaf_17_clock),
    .Q(net108));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2852_ (.D(\u0.cmd[8] ),
    .CLK(clknet_leaf_20_clock),
    .Q(net109));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2853_ (.D(\u0.cmd[9] ),
    .CLK(clknet_leaf_17_clock),
    .Q(net110));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2854_ (.D(\u0.cmd[10] ),
    .CLK(clknet_leaf_19_clock),
    .Q(net96));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2855_ (.D(\u0.cmd[11] ),
    .CLK(clknet_leaf_19_clock),
    .Q(net97));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2856_ (.D(\u0.cmd[12] ),
    .CLK(clknet_leaf_20_clock),
    .Q(net98));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2857_ (.D(\u0.cmd[13] ),
    .CLK(clknet_leaf_19_clock),
    .Q(net99));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2858_ (.D(\u0.cmd[14] ),
    .CLK(clknet_leaf_19_clock),
    .Q(net100));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2859_ (.D(\u0.cmd[15] ),
    .CLK(clknet_leaf_19_clock),
    .Q(net101));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2860_ (.D(\u1.output_active ),
    .CLK(clknet_leaf_7_clock),
    .Q(net192));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2861_ (.D(latch_data),
    .CLK(clknet_leaf_2_clock),
    .Q(\latch_data_sync[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2862_ (.D(\latch_data_sync[0] ),
    .CLK(clknet_leaf_7_clock),
    .Q(\latch_data_sync[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2863_ (.D(control_trigger),
    .CLK(clknet_leaf_15_clock),
    .Q(\control_trigger_sync[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2864_ (.D(\control_trigger_sync[0] ),
    .CLK(clknet_leaf_15_clock),
    .Q(\control_trigger_sync[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2865_ (.D(reset_n),
    .CLK(clknet_leaf_37_clock),
    .Q(\reset_n_sync[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2866_ (.D(\reset_n_sync[0] ),
    .CLK(clknet_leaf_37_clock),
    .Q(\reset_n_sync[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2867_ (.D(_0024_),
    .CLK(clknet_leaf_38_clock),
    .Q(net160));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2868_ (.D(_0025_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u1.col_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2869_ (.D(_0026_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u1.col_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2870_ (.D(_0027_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u1.col_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2871_ (.D(_0028_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u1.col_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2872_ (.D(_0029_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u1.col_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2873_ (.D(_0030_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u1.col_sel[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2874_ (.D(_0031_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u1.col_sel[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2875_ (.D(\u0.latch_cmd ),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.update_cmd ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2876_ (.D(_0022_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u0.write_config_n ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2877_ (.D(_0011_),
    .CLK(clknet_leaf_6_clock),
    .Q(\u0.timer_enable ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2878_ (.D(_0012_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u0.mem_write_n[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2879_ (.D(_0013_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u0.mem_write_n[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2880_ (.D(_0014_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u0.mem_write_n[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2881_ (.D(_0015_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u0.mem_write_n[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2882_ (.D(_0016_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u0.mem_write_n[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2883_ (.D(_0017_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u0.mem_write_n[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2884_ (.D(_0018_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u0.mem_write_n[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2885_ (.D(_0019_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u0.mem_write_n[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2886_ (.D(_0020_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u0.mem_write_n[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2887_ (.D(_0021_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u0.mem_write_n[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2888_ (.D(\u1.ccr1_flag ),
    .CLK(clknet_leaf_17_clock),
    .Q(\u1.u1.impulse_gen[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2889_ (.D(\u1.u1.impulse_gen[0] ),
    .CLK(clknet_leaf_17_clock),
    .Q(\u1.u1.impulse_gen[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2890_ (.D(_0032_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.ccr0[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2891_ (.D(_0033_),
    .CLK(clknet_leaf_25_clock),
    .Q(\u1.ccr0[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2892_ (.D(_0034_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u1.ccr0[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2893_ (.D(_0035_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u1.ccr0[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2894_ (.D(_0036_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.ccr0[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2895_ (.D(_0037_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.ccr0[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2896_ (.D(_0038_),
    .CLK(clknet_leaf_25_clock),
    .Q(\u1.ccr0[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2897_ (.D(_0039_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.ccr0[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2898_ (.D(_0040_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u1.ccr0[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2899_ (.D(_0041_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u1.ccr0[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2900_ (.D(_0042_),
    .CLK(clknet_leaf_25_clock),
    .Q(\u1.ccr0[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2901_ (.D(_0043_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u1.ccr0[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2902_ (.D(_0044_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u1.ccr0[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2903_ (.D(_0045_),
    .CLK(clknet_leaf_28_clock),
    .Q(\u1.ccr0[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2904_ (.D(_0046_),
    .CLK(clknet_leaf_28_clock),
    .Q(\u1.ccr0[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2905_ (.D(_0047_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.ccr0[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2906_ (.D(_0048_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.ccr1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2907_ (.D(_0049_),
    .CLK(clknet_leaf_15_clock),
    .Q(\u1.ccr1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2908_ (.D(_0050_),
    .CLK(clknet_leaf_15_clock),
    .Q(\u1.ccr1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2909_ (.D(_0051_),
    .CLK(clknet_leaf_6_clock),
    .Q(\u1.ccr1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2910_ (.D(_0052_),
    .CLK(clknet_leaf_6_clock),
    .Q(\u1.ccr1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2911_ (.D(_0053_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u1.ccr1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2912_ (.D(_0054_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u1.ccr1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2913_ (.D(_0055_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u1.ccr1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2914_ (.D(_0056_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u1.ccr1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2915_ (.D(_0057_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ccr1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2916_ (.D(_0058_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ccr1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2917_ (.D(_0059_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u1.ccr1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2918_ (.D(_0060_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u1.ccr1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2919_ (.D(_0061_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u1.ccr1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2920_ (.D(_0062_),
    .CLK(clknet_leaf_33_clock),
    .Q(\u1.ccr1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2921_ (.D(_0063_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.ccr1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2922_ (.D(_0064_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u1.ccr1[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2923_ (.D(_0065_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u1.ccr1[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2924_ (.D(_0066_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u1.ccr1[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2925_ (.D(_0067_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u1.ccr1[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2926_ (.D(_0068_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.ccr1[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2927_ (.D(_0069_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.ccr1[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2928_ (.D(_0070_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.ccr1[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2929_ (.D(_0071_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.ccr1[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2930_ (.D(_0072_),
    .CLK(clknet_leaf_25_clock),
    .Q(\u1.ccr1[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2931_ (.D(_0073_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.ccr1[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2932_ (.D(_0074_),
    .CLK(clknet_leaf_25_clock),
    .Q(\u1.ccr1[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2933_ (.D(_0075_),
    .CLK(clknet_leaf_25_clock),
    .Q(\u1.ccr1[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2934_ (.D(_0076_),
    .CLK(clknet_leaf_28_clock),
    .Q(\u1.ccr1[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2935_ (.D(_0077_),
    .CLK(clknet_leaf_28_clock),
    .Q(\u1.ccr1[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2936_ (.D(_0078_),
    .CLK(clknet_leaf_28_clock),
    .Q(\u1.ccr1[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2937_ (.D(_0079_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.ccr1[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2938_ (.D(_0080_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u1.ordering_complete[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2939_ (.D(_0081_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u1.ordering_complete[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2940_ (.D(_0082_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u1.ordering_complete[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2941_ (.D(_0083_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ordering_complete[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2942_ (.D(_0084_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ordering_complete[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2943_ (.D(_0085_),
    .CLK(clknet_leaf_1_clock),
    .Q(\u1.ordering_complete[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2944_ (.D(_0086_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u1.ordering_complete[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2945_ (.D(_0087_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u1.ordering_complete[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2946_ (.D(_0088_),
    .CLK(clknet_leaf_1_clock),
    .Q(\u1.ordering_complete[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2947_ (.D(_0089_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u1.ordering_complete[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2948_ (.D(_0090_),
    .CLK(clknet_leaf_1_clock),
    .Q(\u1.ordering_complete[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2949_ (.D(_0091_),
    .CLK(clknet_leaf_1_clock),
    .Q(\u1.ordering_complete[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2950_ (.D(_0092_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u1.ordering_complete[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2951_ (.D(_0093_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ordering_complete[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2952_ (.D(_0094_),
    .CLK(clknet_leaf_35_clock),
    .Q(\u1.ordering_complete[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2953_ (.D(_0095_),
    .CLK(clknet_leaf_35_clock),
    .Q(\u1.ordering_complete[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2954_ (.D(_0096_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u1.ordering_complete[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2955_ (.D(_0097_),
    .CLK(clknet_leaf_33_clock),
    .Q(\u1.ordering_complete[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2956_ (.D(_0098_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u1.ordering_complete[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2957_ (.D(_0099_),
    .CLK(clknet_leaf_33_clock),
    .Q(\u1.ordering_complete[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2958_ (.D(_0100_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u1.ordering_complete[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2959_ (.D(_0101_),
    .CLK(clknet_leaf_33_clock),
    .Q(\u1.ordering_complete[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2960_ (.D(_0102_),
    .CLK(clknet_leaf_33_clock),
    .Q(\u1.ordering_complete[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2961_ (.D(_0103_),
    .CLK(clknet_leaf_33_clock),
    .Q(\u1.ordering_complete[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2962_ (.D(_0104_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.ordering_complete[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2963_ (.D(_0105_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u1.ordering_complete[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2964_ (.D(_0106_),
    .CLK(clknet_leaf_33_clock),
    .Q(\u1.ordering_complete[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2965_ (.D(_0107_),
    .CLK(clknet_leaf_33_clock),
    .Q(\u1.ordering_complete[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2966_ (.D(_0108_),
    .CLK(clknet_leaf_28_clock),
    .Q(\u1.ordering_complete[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2967_ (.D(_0109_),
    .CLK(clknet_leaf_33_clock),
    .Q(\u1.ordering_complete[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2968_ (.D(_0110_),
    .CLK(clknet_leaf_28_clock),
    .Q(\u1.ordering_complete[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2969_ (.D(_0111_),
    .CLK(clknet_leaf_28_clock),
    .Q(\u1.ordering_complete[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2970_ (.D(_0112_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.row_limit[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2971_ (.D(_0113_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.row_limit[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2972_ (.D(_0114_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.row_limit[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2973_ (.D(_0115_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.row_limit[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2974_ (.D(_0116_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.row_limit[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2975_ (.D(_0117_),
    .CLK(clknet_leaf_15_clock),
    .Q(\u1.row_limit[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2976_ (.D(_0118_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.row_limit[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2977_ (.D(_0119_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u1.col_limit[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2978_ (.D(_0120_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u1.col_limit[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2979_ (.D(_0121_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u1.col_limit[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2980_ (.D(_0122_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u1.col_limit[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2981_ (.D(_0123_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.col_limit[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2982_ (.D(_0124_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u1.col_limit[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2983_ (.D(_0125_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u1.col_limit[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2984_ (.D(_0126_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u1.inverter_select[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2985_ (.D(_0127_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u1.inverter_select[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2986_ (.D(_0128_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u1.inverter_select[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2987_ (.D(_0129_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u1.inverter_select[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2988_ (.D(_0130_),
    .CLK(clknet_leaf_22_clock),
    .Q(\u1.inverter_select[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2989_ (.D(_0131_),
    .CLK(clknet_leaf_22_clock),
    .Q(\u1.inverter_select[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2990_ (.D(_0132_),
    .CLK(clknet_leaf_22_clock),
    .Q(\u1.inverter_select[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2991_ (.D(_0133_),
    .CLK(clknet_leaf_21_clock),
    .Q(\u1.inverter_select[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2992_ (.D(_0134_),
    .CLK(clknet_leaf_22_clock),
    .Q(\u1.inverter_select[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2993_ (.D(_0135_),
    .CLK(clknet_leaf_22_clock),
    .Q(\u1.inverter_select[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2994_ (.D(_0136_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u1.row_col_select[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2995_ (.D(_0137_),
    .CLK(clknet_leaf_21_clock),
    .Q(\u1.row_col_select[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2996_ (.D(_0138_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u1.row_col_select[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2997_ (.D(_0139_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u1.row_col_select[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2998_ (.D(_0140_),
    .CLK(clknet_leaf_21_clock),
    .Q(\u1.row_col_select[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2999_ (.D(_0141_),
    .CLK(clknet_leaf_22_clock),
    .Q(\u1.row_col_select[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3000_ (.D(_0142_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u1.row_col_select[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3001_ (.D(_0143_),
    .CLK(clknet_leaf_21_clock),
    .Q(\u1.row_col_select[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3002_ (.D(_0144_),
    .CLK(clknet_leaf_22_clock),
    .Q(\u1.row_col_select[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3003_ (.D(_0145_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u1.row_col_select[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3004_ (.D(_0146_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u1.ordering_timer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3005_ (.D(_0147_),
    .CLK(clknet_leaf_35_clock),
    .Q(\u1.ordering_timer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3006_ (.D(_0148_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u1.ordering_timer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3007_ (.D(_0149_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u1.ordering_timer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3008_ (.D(_0150_),
    .CLK(clknet_leaf_1_clock),
    .Q(\u1.ordering_timer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3009_ (.D(_0151_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u1.ordering_timer[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3010_ (.D(_0152_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u1.ordering_timer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3011_ (.D(_0153_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u1.ordering_timer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3012_ (.D(_0154_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u1.ordering_timer[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3013_ (.D(_0155_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u1.ordering_timer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3014_ (.D(_0156_),
    .CLK(clknet_leaf_37_clock),
    .Q(\u1.ordering_timer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3015_ (.D(_0157_),
    .CLK(clknet_leaf_37_clock),
    .Q(\u1.ordering_timer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3016_ (.D(_0158_),
    .CLK(clknet_leaf_37_clock),
    .Q(\u1.ordering_timer[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3017_ (.D(_0159_),
    .CLK(clknet_leaf_37_clock),
    .Q(\u1.ordering_timer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3018_ (.D(_0160_),
    .CLK(clknet_leaf_35_clock),
    .Q(\u1.ordering_timer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3019_ (.D(_0161_),
    .CLK(clknet_leaf_35_clock),
    .Q(\u1.ordering_timer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3020_ (.D(_0162_),
    .CLK(clknet_leaf_35_clock),
    .Q(\u1.ordering_timer[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3021_ (.D(_0163_),
    .CLK(clknet_leaf_35_clock),
    .Q(\u1.ordering_timer[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3022_ (.D(_0164_),
    .CLK(clknet_leaf_35_clock),
    .Q(\u1.ordering_timer[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3023_ (.D(_0165_),
    .CLK(clknet_leaf_36_clock),
    .Q(\u1.ordering_timer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3024_ (.D(_0166_),
    .CLK(clknet_leaf_32_clock),
    .Q(\u1.ordering_timer[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3025_ (.D(_0167_),
    .CLK(clknet_leaf_32_clock),
    .Q(\u1.ordering_timer[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3026_ (.D(_0168_),
    .CLK(clknet_leaf_31_clock),
    .Q(\u1.ordering_timer[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3027_ (.D(_0169_),
    .CLK(clknet_leaf_32_clock),
    .Q(\u1.ordering_timer[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3028_ (.D(_0170_),
    .CLK(clknet_leaf_31_clock),
    .Q(\u1.ordering_timer[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3029_ (.D(_0171_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u1.ordering_timer[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3030_ (.D(_0172_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u1.ordering_timer[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3031_ (.D(_0173_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u1.ordering_timer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3032_ (.D(_0174_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u1.ordering_timer[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3033_ (.D(_0175_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u1.ordering_timer[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3034_ (.D(_0176_),
    .CLK(clknet_leaf_33_clock),
    .Q(\u1.ordering_timer[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3035_ (.D(_0177_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u1.ordering_timer[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3036_ (.D(_0178_),
    .CLK(clknet_leaf_15_clock),
    .Q(\u0.cmd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3037_ (.D(_0179_),
    .CLK(clknet_leaf_15_clock),
    .Q(\u0.cmd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3038_ (.D(_0180_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.cmd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3039_ (.D(_0181_),
    .CLK(clknet_leaf_6_clock),
    .Q(\u0.cmd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3040_ (.D(_0182_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.cmd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3041_ (.D(_0183_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u0.cmd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3042_ (.D(_0184_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u0.cmd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3043_ (.D(_0185_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u0.cmd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3044_ (.D(_0186_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u0.cmd[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3045_ (.D(_0187_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u0.cmd[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3046_ (.D(_0188_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u0.cmd[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3047_ (.D(_0189_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u0.cmd[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3048_ (.D(_0190_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u0.cmd[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3049_ (.D(_0191_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u0.cmd[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3050_ (.D(_0192_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u0.cmd[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3051_ (.D(_0193_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u0.cmd[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3052_ (.D(_0194_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.cmd[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3053_ (.D(_0195_),
    .CLK(clknet_leaf_6_clock),
    .Q(\u0.cmd[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3054_ (.D(_0196_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.cmd[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3055_ (.D(_0197_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.cmd[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3056_ (.D(_0198_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.cmd[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _3057_ (.D(_0199_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.cmd[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3058_ (.D(_0200_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u0.cmd[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3059_ (.D(_0201_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u0.cmd[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3060_ (.D(_0202_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u0.cmd[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3061_ (.D(_0203_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u0.cmd[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3062_ (.D(_0204_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u0.cmd[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3063_ (.D(_0205_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u0.cmd[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3064_ (.D(_0206_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u0.cmd[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3065_ (.D(_0207_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u0.cmd[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3066_ (.D(_0208_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u0.cmd[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3067_ (.D(_0209_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u0.cmd[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3068_ (.D(_0023_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u1.output_active ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3069_ (.D(_0210_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u1.row_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3070_ (.D(_0211_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u1.row_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3071_ (.D(_0212_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u1.row_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3072_ (.D(_0213_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u1.row_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3073_ (.D(_0214_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u1.row_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3074_ (.D(_0215_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u1.row_sel[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3075_ (.D(_0216_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u1.row_sel[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3076_ (.D(_0217_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u0.u11.impulse_gen[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3077_ (.D(_0218_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u0.u11.impulse_gen[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3078_ (.D(_0006_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u0.run_state[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3079_ (.D(_0004_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u0.run_state[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3080_ (.D(_0005_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u0.run_state[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3081_ (.D(_0007_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u0.run_state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3082_ (.D(_0008_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u0.run_state[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3083_ (.D(_0009_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u0.run_state[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3084_ (.D(_0010_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u0.run_state[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3085_ (.D(_0219_),
    .CLK(clknet_leaf_38_clock),
    .Q(net149));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3086_ (.D(_0220_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u1.timer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3087_ (.D(_0221_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u1.timer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3088_ (.D(_0222_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u1.timer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3089_ (.D(_0223_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u1.timer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3090_ (.D(_0224_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u1.timer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3091_ (.D(_0225_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.timer[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3092_ (.D(_0226_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u1.timer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3093_ (.D(_0227_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u1.timer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3094_ (.D(_0228_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u1.timer[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3095_ (.D(_0229_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u1.timer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3096_ (.D(_0230_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u1.timer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3097_ (.D(_0231_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u1.timer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3098_ (.D(_0232_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u1.timer[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3099_ (.D(_0233_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.timer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3100_ (.D(_0234_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.timer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3101_ (.D(_0235_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.timer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3102_ (.D(_0236_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.timer[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3103_ (.D(_0237_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.timer[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3104_ (.D(_0238_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u1.timer[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3105_ (.D(_0239_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u1.timer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3106_ (.D(_0240_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.timer[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3107_ (.D(_0241_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.timer[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3108_ (.D(_0242_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.timer[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3109_ (.D(_0243_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.timer[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3110_ (.D(_0244_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.timer[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3111_ (.D(_0245_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u1.timer[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3112_ (.D(_0246_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.timer[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3113_ (.D(_0247_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u1.timer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3114_ (.D(_0248_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u1.timer[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3115_ (.D(_0249_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u1.timer[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3116_ (.D(_0250_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u1.timer[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3117_ (.D(_0251_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u1.timer[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3118_ (.D(net40),
    .CLK(net72),
    .Q(\spi_data_crossing[0].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3119_ (.D(\spi_data_crossing[0].A ),
    .CLK(clknet_leaf_38_clock),
    .Q(\spi_data_crossing[0].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3120_ (.D(net51),
    .CLK(net72),
    .Q(\spi_data_crossing[1].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3121_ (.D(\spi_data_crossing[1].A ),
    .CLK(clknet_leaf_0_clock),
    .Q(\spi_data_crossing[1].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3122_ (.D(net62),
    .CLK(net72),
    .Q(\spi_data_crossing[2].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3123_ (.D(\spi_data_crossing[2].A ),
    .CLK(clknet_leaf_38_clock),
    .Q(\spi_data_crossing[2].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3124_ (.D(net65),
    .CLK(net72),
    .Q(\spi_data_crossing[3].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3125_ (.D(\spi_data_crossing[3].A ),
    .CLK(clknet_leaf_0_clock),
    .Q(\spi_data_crossing[3].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3126_ (.D(net66),
    .CLK(net72),
    .Q(\spi_data_crossing[4].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3127_ (.D(\spi_data_crossing[4].A ),
    .CLK(clknet_leaf_38_clock),
    .Q(\spi_data_crossing[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3128_ (.D(net67),
    .CLK(net72),
    .Q(\spi_data_crossing[5].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3129_ (.D(\spi_data_crossing[5].A ),
    .CLK(clknet_leaf_0_clock),
    .Q(\spi_data_crossing[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3130_ (.D(net68),
    .CLK(net72),
    .Q(\spi_data_crossing[6].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3131_ (.D(\spi_data_crossing[6].A ),
    .CLK(clknet_leaf_0_clock),
    .Q(\spi_data_crossing[6].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3132_ (.D(net69),
    .CLK(net72),
    .Q(\spi_data_crossing[7].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3133_ (.D(\spi_data_crossing[7].A ),
    .CLK(clknet_leaf_2_clock),
    .Q(\spi_data_crossing[7].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3134_ (.D(net70),
    .CLK(net72),
    .Q(\spi_data_crossing[8].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3135_ (.D(\spi_data_crossing[8].A ),
    .CLK(clknet_leaf_2_clock),
    .Q(\spi_data_crossing[8].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3136_ (.D(net71),
    .CLK(net72),
    .Q(\spi_data_crossing[9].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3137_ (.D(\spi_data_crossing[9].A ),
    .CLK(clknet_leaf_2_clock),
    .Q(\spi_data_crossing[9].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3138_ (.D(net41),
    .CLK(net72),
    .Q(\spi_data_crossing[10].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3139_ (.D(\spi_data_crossing[10].A ),
    .CLK(clknet_leaf_2_clock),
    .Q(\spi_data_crossing[10].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3140_ (.D(net42),
    .CLK(net72),
    .Q(\spi_data_crossing[11].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3141_ (.D(\spi_data_crossing[11].A ),
    .CLK(clknet_leaf_2_clock),
    .Q(\spi_data_crossing[11].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3142_ (.D(net43),
    .CLK(net72),
    .Q(\spi_data_crossing[12].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3143_ (.D(\spi_data_crossing[12].A ),
    .CLK(clknet_leaf_2_clock),
    .Q(\spi_data_crossing[12].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3144_ (.D(net44),
    .CLK(net72),
    .Q(\spi_data_crossing[13].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3145_ (.D(\spi_data_crossing[13].A ),
    .CLK(clknet_leaf_2_clock),
    .Q(\spi_data_crossing[13].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3146_ (.D(net45),
    .CLK(net72),
    .Q(\spi_data_crossing[14].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3147_ (.D(\spi_data_crossing[14].A ),
    .CLK(clknet_leaf_2_clock),
    .Q(\spi_data_crossing[14].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3148_ (.D(net46),
    .CLK(net72),
    .Q(\spi_data_crossing[15].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3149_ (.D(\spi_data_crossing[15].A ),
    .CLK(clknet_leaf_2_clock),
    .Q(\spi_data_crossing[15].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3150_ (.D(net47),
    .CLK(net72),
    .Q(\spi_data_crossing[16].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3151_ (.D(\spi_data_crossing[16].A ),
    .CLK(clknet_leaf_7_clock),
    .Q(\spi_data_crossing[16].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3152_ (.D(net48),
    .CLK(net72),
    .Q(\spi_data_crossing[17].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3153_ (.D(\spi_data_crossing[17].A ),
    .CLK(clknet_leaf_8_clock),
    .Q(\spi_data_crossing[17].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3154_ (.D(net49),
    .CLK(net72),
    .Q(\spi_data_crossing[18].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3155_ (.D(\spi_data_crossing[18].A ),
    .CLK(clknet_leaf_8_clock),
    .Q(\spi_data_crossing[18].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3156_ (.D(net50),
    .CLK(net72),
    .Q(\spi_data_crossing[19].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3157_ (.D(\spi_data_crossing[19].A ),
    .CLK(clknet_leaf_8_clock),
    .Q(\spi_data_crossing[19].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3158_ (.D(net52),
    .CLK(net72),
    .Q(\spi_data_crossing[20].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3159_ (.D(\spi_data_crossing[20].A ),
    .CLK(clknet_leaf_8_clock),
    .Q(\spi_data_crossing[20].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3160_ (.D(net53),
    .CLK(net72),
    .Q(\spi_data_crossing[21].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3161_ (.D(\spi_data_crossing[21].A ),
    .CLK(clknet_leaf_8_clock),
    .Q(\spi_data_crossing[21].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3162_ (.D(net54),
    .CLK(net72),
    .Q(\spi_data_crossing[22].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3163_ (.D(\spi_data_crossing[22].A ),
    .CLK(clknet_leaf_9_clock),
    .Q(\spi_data_crossing[22].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3164_ (.D(net55),
    .CLK(net72),
    .Q(\spi_data_crossing[23].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3165_ (.D(\spi_data_crossing[23].A ),
    .CLK(clknet_leaf_10_clock),
    .Q(\spi_data_crossing[23].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3166_ (.D(net56),
    .CLK(net72),
    .Q(\spi_data_crossing[24].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3167_ (.D(\spi_data_crossing[24].A ),
    .CLK(clknet_leaf_10_clock),
    .Q(\spi_data_crossing[24].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3168_ (.D(net57),
    .CLK(net72),
    .Q(\spi_data_crossing[25].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3169_ (.D(\spi_data_crossing[25].A ),
    .CLK(clknet_leaf_10_clock),
    .Q(\spi_data_crossing[25].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3170_ (.D(net58),
    .CLK(net72),
    .Q(\spi_data_crossing[26].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3171_ (.D(\spi_data_crossing[26].A ),
    .CLK(clknet_leaf_10_clock),
    .Q(\spi_data_crossing[26].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3172_ (.D(net59),
    .CLK(net72),
    .Q(\spi_data_crossing[27].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3173_ (.D(\spi_data_crossing[27].A ),
    .CLK(clknet_leaf_10_clock),
    .Q(\spi_data_crossing[27].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3174_ (.D(net60),
    .CLK(net72),
    .Q(\spi_data_crossing[28].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3175_ (.D(\spi_data_crossing[28].A ),
    .CLK(clknet_leaf_11_clock),
    .Q(\spi_data_crossing[28].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3176_ (.D(net61),
    .CLK(net72),
    .Q(\spi_data_crossing[29].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3177_ (.D(\spi_data_crossing[29].A ),
    .CLK(clknet_leaf_12_clock),
    .Q(\spi_data_crossing[29].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3178_ (.D(net63),
    .CLK(net72),
    .Q(\spi_data_crossing[30].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3179_ (.D(\spi_data_crossing[30].A ),
    .CLK(clknet_leaf_10_clock),
    .Q(\spi_data_crossing[30].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3180_ (.D(net64),
    .CLK(net72),
    .Q(\spi_data_crossing[31].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3181_ (.D(\spi_data_crossing[31].A ),
    .CLK(clknet_leaf_10_clock),
    .Q(\spi_data_crossing[31].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3182_ (.D(_0252_),
    .CLK(clknet_leaf_31_clock),
    .Q(net148));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3183_ (.D(_0253_),
    .CLK(clknet_leaf_32_clock),
    .Q(net146));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3184_ (.D(_0254_),
    .CLK(clknet_leaf_36_clock),
    .Q(net144));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3185_ (.D(_0255_),
    .CLK(clknet_leaf_36_clock),
    .Q(net142));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3186_ (.D(_0256_),
    .CLK(clknet_leaf_36_clock),
    .Q(net140));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3187_ (.D(_0257_),
    .CLK(clknet_leaf_37_clock),
    .Q(net157));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3188_ (.D(_0258_),
    .CLK(clknet_leaf_37_clock),
    .Q(net155));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3189_ (.D(_0259_),
    .CLK(clknet_leaf_37_clock),
    .Q(net153));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3190_ (.D(_0260_),
    .CLK(clknet_leaf_38_clock),
    .Q(net151));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3191_ (.D(_0261_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.ccr0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3192_ (.D(_0262_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.ccr0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3193_ (.D(_0263_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u1.ccr0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3194_ (.D(_0264_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.ccr0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3195_ (.D(_0265_),
    .CLK(clknet_leaf_6_clock),
    .Q(\u1.ccr0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3196_ (.D(_0266_),
    .CLK(clknet_leaf_6_clock),
    .Q(\u1.ccr0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3197_ (.D(_0267_),
    .CLK(clknet_leaf_15_clock),
    .Q(\u1.ccr0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3198_ (.D(_0268_),
    .CLK(clknet_leaf_6_clock),
    .Q(\u1.ccr0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3199_ (.D(_0269_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.ccr0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3200_ (.D(_0270_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.ccr0[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3201_ (.D(_0271_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u1.ccr0[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3202_ (.D(_0272_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u1.ccr0[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3203_ (.D(_0273_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u1.ccr0[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3204_ (.D(_0274_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u1.ccr0[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3205_ (.D(_0275_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.ccr0[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3206_ (.D(_0276_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u1.ccr0[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3207_ (.D(_0277_),
    .CLK(clknet_leaf_38_clock),
    .Q(net159));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3208_ (.D(_0278_),
    .CLK(clknet_leaf_38_clock),
    .Q(net158));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3209_ (.D(_0001_),
    .CLK(clknet_leaf_38_clock),
    .Q(net161));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3210_ (.D(_0279_),
    .CLK(clknet_leaf_36_clock),
    .Q(net137));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3211_ (.D(_0003_),
    .CLK(clknet_leaf_37_clock),
    .Q(reset_n));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3212_ (.D(_0002_),
    .CLK(clknet_leaf_37_clock),
    .Q(latch_data));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3213_ (.D(_0000_),
    .CLK(clknet_leaf_36_clock),
    .Q(control_trigger));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3214_ (.D(\u1.inverter_select[0] ),
    .CLK(clknet_leaf_20_clock),
    .Q(net127));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3215_ (.D(\u1.inverter_select[1] ),
    .CLK(clknet_leaf_20_clock),
    .Q(net128));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3216_ (.D(\u1.inverter_select[2] ),
    .CLK(clknet_leaf_22_clock),
    .Q(net129));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3217_ (.D(\u1.inverter_select[3] ),
    .CLK(clknet_leaf_21_clock),
    .Q(net130));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3218_ (.D(\u1.inverter_select[4] ),
    .CLK(clknet_leaf_21_clock),
    .Q(net131));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3219_ (.D(\u1.inverter_select[5] ),
    .CLK(clknet_leaf_21_clock),
    .Q(net132));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3220_ (.D(\u1.inverter_select[6] ),
    .CLK(clknet_leaf_21_clock),
    .Q(net133));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3221_ (.D(\u1.inverter_select[7] ),
    .CLK(clknet_leaf_21_clock),
    .Q(net134));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3222_ (.D(\u1.inverter_select[8] ),
    .CLK(clknet_leaf_21_clock),
    .Q(net135));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3223_ (.D(\u1.inverter_select[9] ),
    .CLK(clknet_leaf_22_clock),
    .Q(net136));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3224_ (.D(\u1.row_col_select[0] ),
    .CLK(clknet_leaf_21_clock),
    .Q(net194));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3225_ (.D(\u1.row_col_select[1] ),
    .CLK(clknet_leaf_21_clock),
    .Q(net195));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3226_ (.D(\u1.row_col_select[2] ),
    .CLK(clknet_leaf_21_clock),
    .Q(net196));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3227_ (.D(\u1.row_col_select[3] ),
    .CLK(clknet_leaf_21_clock),
    .Q(net197));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3228_ (.D(\u1.row_col_select[4] ),
    .CLK(clknet_leaf_21_clock),
    .Q(net198));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3229_ (.D(\u1.row_col_select[5] ),
    .CLK(clknet_leaf_21_clock),
    .Q(net199));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3230_ (.D(\u1.row_col_select[6] ),
    .CLK(clknet_leaf_22_clock),
    .Q(net200));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3231_ (.D(\u1.row_col_select[7] ),
    .CLK(clknet_leaf_21_clock),
    .Q(net201));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3232_ (.D(\u1.row_col_select[8] ),
    .CLK(clknet_leaf_22_clock),
    .Q(net202));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3233_ (.D(\u1.row_col_select[9] ),
    .CLK(clknet_leaf_22_clock),
    .Q(net203));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3234_ (.D(\u0.cmd[16] ),
    .CLK(clknet_leaf_8_clock),
    .Q(net162));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3235_ (.D(\u0.cmd[17] ),
    .CLK(clknet_leaf_12_clock),
    .Q(net163));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3236_ (.D(\u0.cmd[18] ),
    .CLK(clknet_leaf_9_clock),
    .Q(net164));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3237_ (.D(\u0.cmd[19] ),
    .CLK(clknet_leaf_9_clock),
    .Q(net165));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3238_ (.D(\u0.cmd[20] ),
    .CLK(clknet_leaf_10_clock),
    .Q(net166));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3239_ (.D(\u0.cmd[21] ),
    .CLK(clknet_leaf_9_clock),
    .Q(net167));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3240_ (.D(\u0.cmd[22] ),
    .CLK(clknet_leaf_10_clock),
    .Q(net168));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3241_ (.D(\u0.cmd[23] ),
    .CLK(clknet_leaf_10_clock),
    .Q(net169));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3242_ (.D(\u0.cmd[24] ),
    .CLK(clknet_leaf_11_clock),
    .Q(net170));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3243_ (.D(\u0.cmd[25] ),
    .CLK(clknet_leaf_11_clock),
    .Q(net171));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3244_ (.D(\u0.mem_write_n[0] ),
    .CLK(clknet_leaf_11_clock),
    .Q(net182));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3245_ (.D(\u0.mem_write_n[1] ),
    .CLK(clknet_leaf_11_clock),
    .Q(net183));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3246_ (.D(\u0.mem_write_n[2] ),
    .CLK(clknet_leaf_11_clock),
    .Q(net184));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3247_ (.D(\u0.mem_write_n[3] ),
    .CLK(clknet_leaf_11_clock),
    .Q(net185));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3248_ (.D(\u0.mem_write_n[4] ),
    .CLK(clknet_leaf_13_clock),
    .Q(net186));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3249_ (.D(\u0.mem_write_n[5] ),
    .CLK(clknet_leaf_13_clock),
    .Q(net187));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3250_ (.D(\u0.mem_write_n[6] ),
    .CLK(clknet_leaf_12_clock),
    .Q(net188));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3251_ (.D(\u0.mem_write_n[7] ),
    .CLK(clknet_leaf_12_clock),
    .Q(net189));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3252_ (.D(\u0.mem_write_n[8] ),
    .CLK(clknet_leaf_12_clock),
    .Q(net190));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3253_ (.D(\u0.mem_write_n[9] ),
    .CLK(clknet_leaf_12_clock),
    .Q(net191));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3254_ (.I(clknet_leaf_12_clock),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3255_ (.I(clknet_leaf_12_clock),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3256_ (.I(clknet_leaf_12_clock),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3257_ (.I(clknet_leaf_12_clock),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3258_ (.I(clknet_leaf_12_clock),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3259_ (.I(clknet_leaf_12_clock),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3260_ (.I(clknet_leaf_12_clock),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3261_ (.I(clknet_leaf_12_clock),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3262_ (.I(clknet_leaf_12_clock),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3263_ (.I(clknet_leaf_12_clock),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3264_ (.I(net83),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3265_ (.I(net84),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3266_ (.I(net85),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3267_ (.I(net86),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3268_ (.I(net87),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3269_ (.I(net88),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3270_ (.I(net95),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3271_ (.I(net102),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3272_ (.I(net103),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3273_ (.I(net104),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3274_ (.I(net105),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3275_ (.I(net106),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3276_ (.I(net107),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3277_ (.I(net108),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3278_ (.I(net109),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3279_ (.I(net110),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3280_ (.I(net96),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3281_ (.I(net97),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3282_ (.I(net98),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3283_ (.I(net99),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3284_ (.I(net100),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3285_ (.I(net101),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3286_ (.I(net149),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3287_ (.I(net151),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3288_ (.I(net153),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3289_ (.I(net155),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3290_ (.I(net157),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3291_ (.I(net140),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3292_ (.I(net142),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3293_ (.I(net144),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3294_ (.I(net146),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3295_ (.I(net148),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3296_ (.I(net162),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3297_ (.I(net163),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3298_ (.I(net164),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3299_ (.I(net165),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3300_ (.I(net166),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3301_ (.I(net167),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3302_ (.I(net168),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3303_ (.I(net169),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3304_ (.I(net170),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3305_ (.I(net171),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3306_ (.I(net192),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3307_ (.I(net204),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3308_ (.I(net205),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3309_ (.I(net206),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3310_ (.I(net207),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3311_ (.I(net208),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3312_ (.I(net209),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(io_control_trigger_in),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(io_latch_data_in),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(io_reset_n_in),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(la_data_in[0]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(la_data_in[10]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(la_data_in[11]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(la_data_in[12]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(la_data_in[13]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(la_data_in[14]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(la_data_in[15]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(la_data_in[16]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(la_data_in[17]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(la_data_in[1]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(la_data_in[2]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(la_data_in[3]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(la_data_in[4]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(la_data_in[5]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(la_data_in[6]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(la_data_in[7]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(la_data_in[8]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(la_data_in[9]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(la_oenb[0]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(la_oenb[10]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(la_oenb[11]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(la_oenb[12]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(la_oenb[13]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(la_oenb[14]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(la_oenb[15]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(la_oenb[16]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(la_oenb[17]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(la_oenb[1]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(la_oenb[2]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(la_oenb[3]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(la_oenb[4]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(la_oenb[5]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(la_oenb[6]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(la_oenb[7]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(la_oenb[8]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(la_oenb[9]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(spi_data[0]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(spi_data[10]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(spi_data[11]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input43 (.I(spi_data[12]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input44 (.I(spi_data[13]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input45 (.I(spi_data[14]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input46 (.I(spi_data[15]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input47 (.I(spi_data[16]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input48 (.I(spi_data[17]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input49 (.I(spi_data[18]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input50 (.I(spi_data[19]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input51 (.I(spi_data[1]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input52 (.I(spi_data[20]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input53 (.I(spi_data[21]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input54 (.I(spi_data[22]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input55 (.I(spi_data[23]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input56 (.I(spi_data[24]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input57 (.I(spi_data[25]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input58 (.I(spi_data[26]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input59 (.I(spi_data[27]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input60 (.I(spi_data[28]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input61 (.I(spi_data[29]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input62 (.I(spi_data[2]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input63 (.I(spi_data[30]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input64 (.I(spi_data[31]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input65 (.I(spi_data[3]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input66 (.I(spi_data[4]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input67 (.I(spi_data[5]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input68 (.I(spi_data[6]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input69 (.I(spi_data[7]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input70 (.I(spi_data[8]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input71 (.I(spi_data[9]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input72 (.I(spi_data_clock),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output73 (.I(net73),
    .Z(clock_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output74 (.I(net74),
    .Z(clock_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output75 (.I(net75),
    .Z(clock_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output76 (.I(net76),
    .Z(clock_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output77 (.I(net77),
    .Z(clock_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output78 (.I(net78),
    .Z(clock_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output79 (.I(net79),
    .Z(clock_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output80 (.I(net80),
    .Z(clock_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output81 (.I(net81),
    .Z(clock_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output82 (.I(net82),
    .Z(clock_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output83 (.I(net83),
    .Z(col_select_left[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output84 (.I(net84),
    .Z(col_select_left[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output85 (.I(net85),
    .Z(col_select_left[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output86 (.I(net86),
    .Z(col_select_left[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output87 (.I(net87),
    .Z(col_select_left[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output88 (.I(net88),
    .Z(col_select_left[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output89 (.I(net89),
    .Z(col_select_right[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output90 (.I(net90),
    .Z(col_select_right[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output91 (.I(net91),
    .Z(col_select_right[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output92 (.I(net92),
    .Z(col_select_right[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output93 (.I(net93),
    .Z(col_select_right[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output94 (.I(net94),
    .Z(col_select_right[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output95 (.I(net95),
    .Z(data_out_left[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output96 (.I(net96),
    .Z(data_out_left[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output97 (.I(net97),
    .Z(data_out_left[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output98 (.I(net98),
    .Z(data_out_left[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output99 (.I(net99),
    .Z(data_out_left[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output100 (.I(net100),
    .Z(data_out_left[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output101 (.I(net101),
    .Z(data_out_left[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output102 (.I(net102),
    .Z(data_out_left[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output103 (.I(net103),
    .Z(data_out_left[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output104 (.I(net104),
    .Z(data_out_left[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output105 (.I(net105),
    .Z(data_out_left[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output106 (.I(net106),
    .Z(data_out_left[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output107 (.I(net107),
    .Z(data_out_left[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output108 (.I(net108),
    .Z(data_out_left[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output109 (.I(net109),
    .Z(data_out_left[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output110 (.I(net110),
    .Z(data_out_left[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output111 (.I(net111),
    .Z(data_out_right[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output112 (.I(net112),
    .Z(data_out_right[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output113 (.I(net113),
    .Z(data_out_right[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output114 (.I(net114),
    .Z(data_out_right[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output115 (.I(net115),
    .Z(data_out_right[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output116 (.I(net116),
    .Z(data_out_right[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output117 (.I(net117),
    .Z(data_out_right[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output118 (.I(net118),
    .Z(data_out_right[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output119 (.I(net119),
    .Z(data_out_right[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output120 (.I(net120),
    .Z(data_out_right[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output121 (.I(net121),
    .Z(data_out_right[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output122 (.I(net122),
    .Z(data_out_right[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output123 (.I(net123),
    .Z(data_out_right[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output124 (.I(net124),
    .Z(data_out_right[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output125 (.I(net125),
    .Z(data_out_right[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output126 (.I(net126),
    .Z(data_out_right[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output127 (.I(net127),
    .Z(inverter_select[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output128 (.I(net128),
    .Z(inverter_select[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output129 (.I(net129),
    .Z(inverter_select[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output130 (.I(net130),
    .Z(inverter_select[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output131 (.I(net131),
    .Z(inverter_select[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output132 (.I(net132),
    .Z(inverter_select[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output133 (.I(net133),
    .Z(inverter_select[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output134 (.I(net134),
    .Z(inverter_select[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output135 (.I(net135),
    .Z(inverter_select[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output136 (.I(net136),
    .Z(inverter_select[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output137 (.I(net137),
    .Z(io_control_trigger_oeb));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output138 (.I(net138),
    .Z(io_driver_io_oeb[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output139 (.I(net139),
    .Z(io_driver_io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output140 (.I(net140),
    .Z(io_driver_io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output141 (.I(net141),
    .Z(io_driver_io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output142 (.I(net142),
    .Z(io_driver_io_oeb[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output143 (.I(net143),
    .Z(io_driver_io_oeb[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output144 (.I(net144),
    .Z(io_driver_io_oeb[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output145 (.I(net145),
    .Z(io_driver_io_oeb[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output146 (.I(net146),
    .Z(io_driver_io_oeb[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output147 (.I(net147),
    .Z(io_driver_io_oeb[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output148 (.I(net148),
    .Z(io_driver_io_oeb[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output149 (.I(net149),
    .Z(io_driver_io_oeb[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output150 (.I(net150),
    .Z(io_driver_io_oeb[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output151 (.I(net151),
    .Z(io_driver_io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output152 (.I(net152),
    .Z(io_driver_io_oeb[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output153 (.I(net153),
    .Z(io_driver_io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output154 (.I(net154),
    .Z(io_driver_io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output155 (.I(net155),
    .Z(io_driver_io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output156 (.I(net156),
    .Z(io_driver_io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output157 (.I(net157),
    .Z(io_driver_io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output158 (.I(net158),
    .Z(io_latch_data_oeb));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output159 (.I(net159),
    .Z(io_reset_n_oeb));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output160 (.I(net160),
    .Z(io_update_cycle_complete_oeb));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output161 (.I(net161),
    .Z(io_update_cycle_complete_out));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output162 (.I(net162),
    .Z(mem_address_left[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output163 (.I(net163),
    .Z(mem_address_left[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output164 (.I(net164),
    .Z(mem_address_left[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output165 (.I(net165),
    .Z(mem_address_left[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output166 (.I(net166),
    .Z(mem_address_left[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output167 (.I(net167),
    .Z(mem_address_left[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output168 (.I(net168),
    .Z(mem_address_left[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output169 (.I(net169),
    .Z(mem_address_left[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output170 (.I(net170),
    .Z(mem_address_left[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output171 (.I(net171),
    .Z(mem_address_left[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output172 (.I(net172),
    .Z(mem_address_right[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output173 (.I(net173),
    .Z(mem_address_right[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output174 (.I(net174),
    .Z(mem_address_right[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output175 (.I(net175),
    .Z(mem_address_right[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output176 (.I(net176),
    .Z(mem_address_right[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output177 (.I(net177),
    .Z(mem_address_right[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output178 (.I(net178),
    .Z(mem_address_right[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output179 (.I(net179),
    .Z(mem_address_right[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output180 (.I(net180),
    .Z(mem_address_right[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output181 (.I(net181),
    .Z(mem_address_right[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output182 (.I(net182),
    .Z(mem_write_n[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output183 (.I(net183),
    .Z(mem_write_n[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output184 (.I(net184),
    .Z(mem_write_n[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output185 (.I(net185),
    .Z(mem_write_n[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output186 (.I(net186),
    .Z(mem_write_n[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output187 (.I(net187),
    .Z(mem_write_n[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output188 (.I(net188),
    .Z(mem_write_n[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output189 (.I(net189),
    .Z(mem_write_n[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output190 (.I(net190),
    .Z(mem_write_n[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output191 (.I(net191),
    .Z(mem_write_n[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output192 (.I(net192),
    .Z(output_active_left));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output193 (.I(net193),
    .Z(output_active_right));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output194 (.I(net194),
    .Z(row_col_select[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output195 (.I(net195),
    .Z(row_col_select[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output196 (.I(net196),
    .Z(row_col_select[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output197 (.I(net197),
    .Z(row_col_select[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output198 (.I(net198),
    .Z(row_col_select[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output199 (.I(net199),
    .Z(row_col_select[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output200 (.I(net200),
    .Z(row_col_select[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output201 (.I(net201),
    .Z(row_col_select[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output202 (.I(net202),
    .Z(row_col_select[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output203 (.I(net203),
    .Z(row_col_select[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output204 (.I(net204),
    .Z(row_select_left[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output205 (.I(net205),
    .Z(row_select_left[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output206 (.I(net206),
    .Z(row_select_left[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output207 (.I(net207),
    .Z(row_select_left[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output208 (.I(net208),
    .Z(row_select_left[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output209 (.I(net209),
    .Z(row_select_left[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output210 (.I(net210),
    .Z(row_select_right[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output211 (.I(net211),
    .Z(row_select_right[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output212 (.I(net212),
    .Z(row_select_right[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output213 (.I(net213),
    .Z(row_select_right[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output214 (.I(net214),
    .Z(row_select_right[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output215 (.I(net215),
    .Z(row_select_right[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_clock (.I(clknet_2_1__leaf_clock),
    .Z(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_clock (.I(clknet_2_2__leaf_clock),
    .Z(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_clock (.I(clknet_2_3__leaf_clock),
    .Z(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_clock (.I(clknet_2_2__leaf_clock),
    .Z(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_clock (.I(clknet_2_2__leaf_clock),
    .Z(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_clock (.I(clknet_2_2__leaf_clock),
    .Z(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_clock (.I(clknet_2_2__leaf_clock),
    .Z(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_clock (.I(clknet_2_2__leaf_clock),
    .Z(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_clock (.I(clknet_2_2__leaf_clock),
    .Z(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_clock (.I(clknet_2_2__leaf_clock),
    .Z(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_clock (.I(clknet_2_0__leaf_clock),
    .Z(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clock (.I(clock),
    .Z(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_clock (.I(clknet_0_clock),
    .Z(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_clock (.I(clknet_0_clock),
    .Z(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_clock (.I(clknet_0_clock),
    .Z(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_clock (.I(clknet_0_clock),
    .Z(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__D (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__D (.I(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__D (.I(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__D (.I(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__D (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__D (.I(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__D (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__D (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__D (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__D (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__D (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__D (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__D (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3182__D (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__D (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3184__D (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__D (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__D (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__D (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__D (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__D (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3190__D (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A3 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__A3 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__A2 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__A1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__B (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__A3 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__A1 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__B2 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__A1 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__A4 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A2 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A4 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__I (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1812__I (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__A3 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1831__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1828__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1839__A3 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__A1 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__A2 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A3 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__A1 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1828__A2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A4 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A3 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__A2 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__A1 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__A1 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1849__A1 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1859__B2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1857__A2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1859__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__C (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__A1 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A1 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__B (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1880__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__I (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__I1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1955__I1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__I1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1904__I (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__I (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1939__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1920__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1898__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__S (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__S (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__S (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__S (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__I1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__I1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__I1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__I1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__I (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1930__S (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1927__S (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1905__I (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1925__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1922__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2794__I1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__I0 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__I1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1908__A1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1947__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1911__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1908__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__I1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__I0 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__I0 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1911__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__I0 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__I0 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__I1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__I1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2213__I0 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__I0 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__I1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__I1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__I0 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A1 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A1 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__A1 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__A1 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__I1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__I0 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__I1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1927__I1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__I1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__I0 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__I1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1930__I1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__A2 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__A2 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__A2 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1935__A2 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__I1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1934__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1937__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__B (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__I0 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2033__I1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__I1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A1 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__I1 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1996__A1 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__A1 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__I (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1972__I (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__I (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1954__I (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1996__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__S (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1955__S (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__S (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1964__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__A1 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__A1 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__I (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__A1 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__I (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__B (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__I (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__I (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__A2 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__A2 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__A2 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A2 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__I (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2004__I (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1999__I (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__S (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__S (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__S (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2023__I (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__I (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__I (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__S (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__S (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__S (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__S (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__A1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__A1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__A1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2027__A2 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__A2 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__A2 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__A2 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2029__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__B (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__B (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__S (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2033__S (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__S (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__S (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__I0 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__I0 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__I1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__I (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__I (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__I (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2044__I (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__A2 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__A2 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A2 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__A2 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__I (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2090__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A1 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__I0 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__I0 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2055__I0 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2064__S (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__S (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__S (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2055__S (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__I0 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__I0 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__I0 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__I0 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__I0 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__I0 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__I0 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__I0 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2064__I0 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2067__I (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__A1 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__I0 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__I0 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__I0 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__S (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__S (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__S (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__S (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__A1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__I0 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__I0 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__I0 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__I0 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__I0 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__I0 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__I0 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__I0 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__I0 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2083__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2081__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__I (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__I (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__S (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__S (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__I (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__I (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2107__A2 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2105__A2 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__A2 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__A2 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2134__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__S (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__S (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__S (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__S (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2132__A2 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__A2 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__A2 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__A2 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__B2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__A1 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2131__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__A1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__I0 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__I0 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2140__I0 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__I (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__S (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__S (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__I (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__I0 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__I0 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2143__I0 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2162__I (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2160__I (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__S (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__S (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__S (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__I (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__B (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__B (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__S (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__S (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2178__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__S (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__S (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__I (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__I (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__S (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__S (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2213__S (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__S (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__B2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__B (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A2 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A3 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A3 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2252__B (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2252__C (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__A2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2278__A2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2268__A2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__I (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__I (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__I (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__B (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__B (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__B1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__B1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2278__B1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2268__B1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__B (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__S (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__S (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__S (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__I (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__I (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__I (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__I (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__I (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2390__I (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__I (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2287__I (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__I (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__I (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__I (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__I (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__A4 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__A3 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__I (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__I (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__I (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__I (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__I (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__I (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2329__I (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__I (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__I (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__A1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__A1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__A1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__B1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__B1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__B1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__B1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__A3 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A2 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__I (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A3 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__A2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__A2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2358__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__B1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__B1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__B1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__B1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__A4 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__A4 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2398__A3 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__I (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A3 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__B (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__B2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__B (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__I (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A2 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__S (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__S (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__S (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__C (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__C (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__A3 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__I (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A3 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__B (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__C (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__I (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A2 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__C (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__B1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__B1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__B1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__B1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__A2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__A2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__A4 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__I (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A4 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2429__I (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A3 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__A2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__B (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__A1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__B1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__B1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__B1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__B1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A2 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__A3 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A3 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__A3 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A3 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__A3 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A4 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__A3 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A4 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A4 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A2 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__I (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__B (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__A2 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A2 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A3 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__B1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A3 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A2 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__I (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__I (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__I (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__I (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__I (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__I (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__I (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__I (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__I (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__A2 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A2 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__A2 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A2 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__B1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__B1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__B1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__B1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__B1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__B1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__B1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__B1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A2 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__A2 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__A1 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A1 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A1 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A1 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__I (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2640__B (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__B (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__B (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A2 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__A2 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__B2 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__B (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__B2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__A3 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__I (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__I (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__I (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__I (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__C (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__C (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__C (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2667__I (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__A1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__A1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__A1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__A2 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A3 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__A2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__A2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__A3 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__A1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__I (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__I (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2700__I (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__I (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A4 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__A3 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__I (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__A2 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A2 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__A2 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2703__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__A4 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__A2 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__A2 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__A2 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__A4 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__A3 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__A3 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__A3 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__A4 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__A2 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__A3 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__A3 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__C (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__C (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__C (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__I (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__I (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__I (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__I (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__S (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__S (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__S (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__I (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2823__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2821__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A2 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__A2 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A2 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__A2 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2817__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2814__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2821__B (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2827__I (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2829__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__I (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1417__I (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A4 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1533__A3 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1418__A3 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1544__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1530__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1525__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1522__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1527__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1420__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1428__A1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1423__B1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__I (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__B1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__B2 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1437__B2 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1444__B2 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1437__A2 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__A1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__C (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1444__B1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__A1 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1519__A1 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1458__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1449__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2132__A1 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1455__B2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1458__B1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1470__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A3 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A1 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__I (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1465__A1 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1464__B1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A3 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2252__A1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__A2 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1519__A2 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2398__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2376__I (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__I (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1474__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__A1 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__A2 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1480__B2 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__B (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1495__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2331__A1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__A1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1492__B1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1490__A1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__I1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1490__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__A1 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__B1 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1493__A1 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1490__B1 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__I1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1493__A2 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1490__B2 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1519__A3 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1505__B1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__B1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__B (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1502__A2 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1512__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1505__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__B2 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1505__C (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A2 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1507__A3 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1518__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__B (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1518__A3 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1514__I (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1786__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1543__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1520__I (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__B1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1528__A2 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A3 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__A3 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1534__B (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A2 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__A2 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__B2 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__A2 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1546__I (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1566__B2 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1548__I (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1554__B2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__A2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1567__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1554__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1566__A2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__B2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1563__A2 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1569__A3 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A3 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1568__A1 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__A2 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__A1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__A2 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__B2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__B2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__B1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1979__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__B1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__C (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1604__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A3 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__B2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1587__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__I (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__B (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1603__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1598__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A3 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__I (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1598__A2 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A2 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1603__A2 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__B (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__A1 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__A1 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__A1 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__B2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__B1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1628__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A2 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1620__A2 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__B2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1620__B2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1984__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1657__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1633__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1981__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1633__B1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__B (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__B2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1637__B2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__A1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1647__A1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__B1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1659__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__B2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__B2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__B2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__B2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__A2 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2640__A1 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__B (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__I (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__B (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__A2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__B2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__A1 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__A1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__A3 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1671__A1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__B2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__A1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__B (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2814__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__A2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__B (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__B1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__A2 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1699__A2 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__B2 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1699__A3 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1696__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__B1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__B (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1705__I (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__B2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__A2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__I (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1714__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1773__B (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__A3 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__A1 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1773__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__A3 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__B1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1757__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1935__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__B1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1729__B1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__A2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__I (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__B2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1729__B2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__C (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__A1 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A2 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1947__A1 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__B1 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1759__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1754__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__B2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__B (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1769__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__B2 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__A1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__B (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__A1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__A1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__B (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__I (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__I (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1786__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__A1 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1792__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A2 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clock_I (.I(clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__D (.I(control_trigger));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1523__A2 (.I(control_trigger));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1419__A2 (.I(control_trigger));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_control_trigger_in));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_latch_data_in));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_reset_n_in));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(la_data_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(la_data_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(la_data_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(la_data_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(la_data_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(la_data_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(la_data_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(la_data_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(la_data_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(la_data_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(la_data_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(la_data_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(la_data_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(la_data_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(la_data_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(la_data_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(la_data_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(la_data_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(la_oenb[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(la_oenb[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(la_oenb[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(la_oenb[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(la_oenb[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(la_oenb[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(la_oenb[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(la_oenb[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(la_oenb[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(la_oenb[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(la_oenb[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(la_oenb[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(la_oenb[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(la_oenb[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(la_oenb[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(la_oenb[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(la_oenb[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(la_oenb[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__D (.I(latch_data));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A2 (.I(latch_data));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(spi_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(spi_data[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(spi_data[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(spi_data[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(spi_data[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(spi_data[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(spi_data[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(spi_data[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(spi_data[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(spi_data[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(spi_data[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(spi_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(spi_data[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(spi_data[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(spi_data[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(spi_data[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(spi_data[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(spi_data[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(spi_data[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(spi_data[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(spi_data[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(spi_data[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(spi_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(spi_data[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(spi_data[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(spi_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(spi_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(spi_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(spi_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(spi_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(spi_data[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(spi_data[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(spi_data_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__B2 (.I(\spi_data_crossing[0].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__D (.I(\spi_data_crossing[10].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__B2 (.I(\spi_data_crossing[11].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__B2 (.I(\spi_data_crossing[12].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__B2 (.I(\spi_data_crossing[13].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__B2 (.I(\spi_data_crossing[14].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__B2 (.I(\spi_data_crossing[15].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__B2 (.I(\spi_data_crossing[16].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__B2 (.I(\spi_data_crossing[17].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__B2 (.I(\spi_data_crossing[19].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__D (.I(\spi_data_crossing[1].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__B2 (.I(\spi_data_crossing[1].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__B2 (.I(\spi_data_crossing[21].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__B2 (.I(\spi_data_crossing[24].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__D (.I(\spi_data_crossing[25].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__D (.I(\spi_data_crossing[26].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__B2 (.I(\spi_data_crossing[26].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__D (.I(\spi_data_crossing[27].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__D (.I(\spi_data_crossing[28].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__D (.I(\spi_data_crossing[29].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__B2 (.I(\spi_data_crossing[2].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__B2 (.I(\spi_data_crossing[30].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__B2 (.I(\spi_data_crossing[31].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__D (.I(\spi_data_crossing[3].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__B2 (.I(\spi_data_crossing[3].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__B2 (.I(\spi_data_crossing[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__B2 (.I(\spi_data_crossing[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__B2 (.I(\spi_data_crossing[6].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__B2 (.I(\spi_data_crossing[7].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__D (.I(\spi_data_crossing[9].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__D (.I(\u0.cmd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__I (.I(\u0.cmd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1889__I (.I(\u0.cmd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__D (.I(\u0.cmd[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__A1 (.I(\u0.cmd[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__A1 (.I(\u0.cmd[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2081__A1 (.I(\u0.cmd[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1933__I (.I(\u0.cmd[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__D (.I(\u0.cmd[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__A1 (.I(\u0.cmd[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__A1 (.I(\u0.cmd[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2083__A1 (.I(\u0.cmd[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1936__I (.I(\u0.cmd[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__D (.I(\u0.cmd[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__A1 (.I(\u0.cmd[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__I (.I(\u0.cmd[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__A1 (.I(\u0.cmd[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__A1 (.I(\u0.cmd[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__D (.I(\u0.cmd[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A1 (.I(\u0.cmd[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2131__A1 (.I(\u0.cmd[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__A1 (.I(\u0.cmd[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1942__I (.I(\u0.cmd[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__D (.I(\u0.cmd[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__A1 (.I(\u0.cmd[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__A1 (.I(\u0.cmd[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__A1 (.I(\u0.cmd[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1945__I (.I(\u0.cmd[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2859__D (.I(\u0.cmd[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__A1 (.I(\u0.cmd[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__A1 (.I(\u0.cmd[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__A1 (.I(\u0.cmd[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__I (.I(\u0.cmd[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__D (.I(\u0.cmd[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2039__I (.I(\u0.cmd[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__A1 (.I(\u0.cmd[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1890__I (.I(\u0.cmd[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3235__D (.I(\u0.cmd[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__I (.I(\u0.cmd[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__I (.I(\u0.cmd[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__D (.I(\u0.cmd[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__A1 (.I(\u0.cmd[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__A1 (.I(\u0.cmd[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__A2 (.I(\u0.cmd[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__D (.I(\u0.cmd[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__A1 (.I(\u0.cmd[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__A1 (.I(\u0.cmd[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__A1 (.I(\u0.cmd[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__I (.I(\u0.cmd[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__D (.I(\u0.cmd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__I (.I(\u0.cmd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__I (.I(\u0.cmd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__D (.I(\u0.cmd[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A1 (.I(\u0.cmd[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__A3 (.I(\u0.cmd[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__A4 (.I(\u0.cmd[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__D (.I(\u0.cmd[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__A1 (.I(\u0.cmd[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__A2 (.I(\u0.cmd[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__A3 (.I(\u0.cmd[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__A2 (.I(\u0.cmd[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1821__A2 (.I(\u0.cmd[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__A1 (.I(\u0.cmd[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1531__I (.I(\u0.cmd[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__D (.I(\u0.cmd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1961__I (.I(\u0.cmd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1906__I (.I(\u0.cmd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A1 (.I(\u0.cmd[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__I (.I(\u0.cmd[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1533__A2 (.I(\u0.cmd[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1418__A2 (.I(\u0.cmd[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__D (.I(\u0.cmd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__I (.I(\u0.cmd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__I (.I(\u0.cmd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__D (.I(\u0.cmd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__I (.I(\u0.cmd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__I (.I(\u0.cmd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__D (.I(\u0.cmd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__I (.I(\u0.cmd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1916__I (.I(\u0.cmd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__D (.I(\u0.cmd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__I (.I(\u0.cmd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1919__I (.I(\u0.cmd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2851__D (.I(\u0.cmd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__A1 (.I(\u0.cmd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__I (.I(\u0.cmd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__I (.I(\u0.cmd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__D (.I(\u0.cmd[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__I (.I(\u0.cmd[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__A1 (.I(\u0.cmd[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__I (.I(\u0.cmd[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__D (.I(\u0.cmd[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__I (.I(\u0.cmd[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A1 (.I(\u0.cmd[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1929__I (.I(\u0.cmd[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__D (.I(\u0.latch_cmd ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__A2 (.I(\u0.latch_cmd ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__A2 (.I(\u0.latch_cmd ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1785__I (.I(\u0.timer_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1594__I (.I(\u0.timer_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__I (.I(\u1.ccr0[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__B1 (.I(\u1.ccr0[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__I (.I(\u1.ccr0[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1680__A2 (.I(\u1.ccr0[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__A2 (.I(\u1.ccr0[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1927__I0 (.I(\u1.ccr0[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__B1 (.I(\u1.ccr0[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1730__B1 (.I(\u1.ccr0[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1930__I0 (.I(\u1.ccr0[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__B1 (.I(\u1.ccr0[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1730__A2 (.I(\u1.ccr0[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2794__I0 (.I(\u1.ccr0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A2 (.I(\u1.ccr0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__B1 (.I(\u1.ccr0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__A2 (.I(\u1.ccr0[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__A2 (.I(\u1.ccr0[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__I (.I(\u1.ccr0[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__I0 (.I(\u1.ccr0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__A2 (.I(\u1.ccr0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__A2 (.I(\u1.ccr0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__I (.I(\u1.ccr0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__A2 (.I(\u1.ccr0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__I0 (.I(\u1.ccr0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__A2 (.I(\u1.ccr0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__B1 (.I(\u1.ccr0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__I0 (.I(\u1.ccr0[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__A2 (.I(\u1.ccr0[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__A2 (.I(\u1.ccr0[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__B1 (.I(\u1.ccr1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__I0 (.I(\u1.ccr1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A1 (.I(\u1.ccr1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__B1 (.I(\u1.ccr1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__I (.I(\u1.ccr1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__C1 (.I(\u1.ccr1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__I0 (.I(\u1.ccr1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__A1 (.I(\u1.ccr1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1592__B1 (.I(\u1.ccr1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__A1 (.I(\u1.ccr1[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__I0 (.I(\u1.ccr1[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__A1 (.I(\u1.ccr1[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1552__A1 (.I(\u1.ccr1[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A1 (.I(\u1.ccr1[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__I0 (.I(\u1.ccr1[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1566__A1 (.I(\u1.ccr1[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__B1 (.I(\u1.ccr1[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2033__I0 (.I(\u1.ccr1[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__A1 (.I(\u1.ccr1[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__B1 (.I(\u1.ccr1[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__I0 (.I(\u1.ccr1[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1554__B1 (.I(\u1.ccr1[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__A1 (.I(\u1.ccr1[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__I0 (.I(\u1.ccr1[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1567__A1 (.I(\u1.ccr1[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1554__A1 (.I(\u1.ccr1[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1582__I (.I(\u1.ccr1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1574__A1 (.I(\u1.ccr1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__A1 (.I(\u1.ccr1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1581__I (.I(\u1.ccr1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__A1 (.I(\u1.ccr1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A1 (.I(\u1.ccr1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1631__I (.I(\u1.ccr1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__I1 (.I(\u1.col_limit[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__B2 (.I(\u1.col_limit[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__B2 (.I(\u1.col_limit[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__I1 (.I(\u1.col_limit[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__A2 (.I(\u1.col_limit[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1849__A2 (.I(\u1.col_limit[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__D (.I(\u1.col_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1859__B1 (.I(\u1.col_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1854__I (.I(\u1.col_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__D (.I(\u1.col_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__B (.I(\u1.col_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__A2 (.I(\u1.col_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1857__B1 (.I(\u1.col_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1853__I (.I(\u1.col_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2842__D (.I(\u1.col_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__A1 (.I(\u1.col_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1881__A1 (.I(\u1.col_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1851__I (.I(\u1.col_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__D (.I(\u1.inverter_select[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__I1 (.I(\u1.inverter_select[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__D (.I(\u1.inverter_select[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__I1 (.I(\u1.inverter_select[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__D (.I(\u1.inverter_select[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__I1 (.I(\u1.inverter_select[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2358__A1 (.I(\u1.ordering_complete[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__I1 (.I(\u1.ordering_complete[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1482__A2 (.I(\u1.ordering_complete[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1481__B2 (.I(\u1.ordering_complete[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__I0 (.I(\u1.ordering_complete[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__I1 (.I(\u1.ordering_complete[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1481__A2 (.I(\u1.ordering_complete[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1477__B2 (.I(\u1.ordering_complete[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__I0 (.I(\u1.ordering_complete[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A2 (.I(\u1.ordering_complete[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1472__I (.I(\u1.ordering_complete[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A1 (.I(\u1.ordering_complete[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__I1 (.I(\u1.ordering_complete[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1431__A2 (.I(\u1.ordering_complete[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1426__B2 (.I(\u1.ordering_complete[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__I0 (.I(\u1.ordering_complete[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__I1 (.I(\u1.ordering_complete[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1428__B2 (.I(\u1.ordering_complete[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1426__A2 (.I(\u1.ordering_complete[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__A1 (.I(\u1.ordering_complete[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__I1 (.I(\u1.ordering_complete[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1428__A2 (.I(\u1.ordering_complete[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1423__B2 (.I(\u1.ordering_complete[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A1 (.I(\u1.ordering_complete[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__I1 (.I(\u1.ordering_complete[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1461__I (.I(\u1.ordering_complete[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__I0 (.I(\u1.ordering_complete[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__I1 (.I(\u1.ordering_complete[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__A2 (.I(\u1.ordering_complete[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1464__B2 (.I(\u1.ordering_complete[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A1 (.I(\u1.ordering_complete[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__I (.I(\u1.ordering_complete[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__B2 (.I(\u1.ordering_complete[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1464__A2 (.I(\u1.ordering_complete[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__I (.I(\u1.ordering_complete[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__A2 (.I(\u1.ordering_complete[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1450__B2 (.I(\u1.ordering_complete[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A1 (.I(\u1.ordering_complete[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__I1 (.I(\u1.ordering_complete[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1452__B2 (.I(\u1.ordering_complete[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1450__A2 (.I(\u1.ordering_complete[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__A1 (.I(\u1.ordering_complete[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1454__I (.I(\u1.ordering_complete[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1452__A2 (.I(\u1.ordering_complete[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__A1 (.I(\u1.ordering_complete[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__I1 (.I(\u1.ordering_complete[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1512__A2 (.I(\u1.ordering_complete[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1505__A2 (.I(\u1.ordering_complete[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__A1 (.I(\u1.ordering_complete[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__I1 (.I(\u1.ordering_complete[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1506__A2 (.I(\u1.ordering_complete[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1501__B2 (.I(\u1.ordering_complete[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__B2 (.I(\u1.ordering_complete[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1487__I (.I(\u1.ordering_complete[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1492__B2 (.I(\u1.ordering_complete[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1485__I (.I(\u1.ordering_complete[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A1 (.I(\u1.ordering_timer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1513__I (.I(\u1.ordering_timer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1510__A1 (.I(\u1.ordering_timer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__I (.I(\u1.ordering_timer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__A1 (.I(\u1.ordering_timer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1480__B1 (.I(\u1.ordering_timer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2398__A2 (.I(\u1.ordering_timer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__I (.I(\u1.ordering_timer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1475__I (.I(\u1.ordering_timer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1474__B1 (.I(\u1.ordering_timer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1480__A1 (.I(\u1.ordering_timer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1471__I (.I(\u1.ordering_timer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A2 (.I(\u1.ordering_timer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__I (.I(\u1.ordering_timer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1515__A1 (.I(\u1.ordering_timer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1510__B1 (.I(\u1.ordering_timer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__I (.I(\u1.ordering_timer[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__B1 (.I(\u1.ordering_timer[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1462__I (.I(\u1.ordering_timer[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A1 (.I(\u1.ordering_timer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A1 (.I(\u1.ordering_timer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__A1 (.I(\u1.ordering_timer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1447__I (.I(\u1.ordering_timer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A1 (.I(\u1.ordering_timer[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A1 (.I(\u1.ordering_timer[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1446__I (.I(\u1.ordering_timer[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A2 (.I(\u1.ordering_timer[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__B (.I(\u1.ordering_timer[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1455__B1 (.I(\u1.ordering_timer[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1451__I (.I(\u1.ordering_timer[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__I (.I(\u1.ordering_timer[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1458__A1 (.I(\u1.ordering_timer[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1449__A1 (.I(\u1.ordering_timer[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__A1 (.I(\u1.ordering_timer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A1 (.I(\u1.ordering_timer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A1 (.I(\u1.ordering_timer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1500__I (.I(\u1.ordering_timer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__D (.I(\u1.row_col_select[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__I1 (.I(\u1.row_col_select[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__D (.I(\u1.row_col_select[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__I1 (.I(\u1.row_col_select[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__D (.I(\u1.row_col_select[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__I1 (.I(\u1.row_col_select[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__D (.I(\u1.row_col_select[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__I1 (.I(\u1.row_col_select[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__B1 (.I(\u1.row_limit[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__A1 (.I(\u1.row_limit[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__I1 (.I(\u1.row_limit[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__B1 (.I(\u1.row_limit[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__A1 (.I(\u1.row_limit[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__I1 (.I(\u1.row_limit[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__D (.I(\u1.row_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A1 (.I(\u1.row_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__A1 (.I(\u1.row_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__I (.I(\u1.row_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__D (.I(\u1.row_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__A1 (.I(\u1.row_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A1 (.I(\u1.row_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__B2 (.I(\u1.row_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__I (.I(\u1.row_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1683__I (.I(\u1.timer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__A2 (.I(\u1.timer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1640__I (.I(\u1.timer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1686__I (.I(\u1.timer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1638__I (.I(\u1.timer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1637__A2 (.I(\u1.timer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__A2 (.I(\u1.timer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__I (.I(\u1.timer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1621__A2 (.I(\u1.timer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__I (.I(\u1.timer[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__B2 (.I(\u1.timer[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1611__I (.I(\u1.timer[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1609__B2 (.I(\u1.timer[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__A1 (.I(\u1.timer[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__B (.I(\u1.timer[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__A4 (.I(\u1.timer[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1547__I (.I(\u1.timer[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__I (.I(\u1.timer[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1545__I (.I(\u1.timer[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1728__I (.I(\u1.timer[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__I (.I(\u1.timer[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1561__B2 (.I(\u1.timer[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1561__A2 (.I(\u1.timer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__I (.I(\u1.timer[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1796__I (.I(\u1.timer[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1742__B2 (.I(\u1.timer[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1555__I (.I(\u1.timer[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__I (.I(\u1.timer[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A3 (.I(\u1.timer[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1742__A1 (.I(\u1.timer[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1550__I (.I(\u1.timer[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A1 (.I(\u1.timer[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A2 (.I(\u1.timer[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__B2 (.I(\u1.timer[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1549__I (.I(\u1.timer[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A2 (.I(\u1.timer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1670__I (.I(\u1.timer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__B2 (.I(\u1.timer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__I (.I(\u1.timer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A1 (.I(\u1.timer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__I (.I(\u1.timer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__A2 (.I(\u1.timer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1575__I (.I(\u1.timer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__I1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__I1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2826__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2830__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__I0 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__I0 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__I0 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__S (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__S (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3178__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3176__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3174__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3172__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3170__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3168__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3164__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3162__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3158__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3156__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3154__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3150__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3146__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3144__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3142__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3138__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3136__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3134__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3130__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3126__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3124__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3118__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output87_I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3268__I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output88_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3269__I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output91_I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output95_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3270__I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output96_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3280__I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output97_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3281__I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output98_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output99_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output100_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output101_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3285__I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output102_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3271__I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output103_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output104_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3273__I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output105_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3274__I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output106_I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output107_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output108_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output109_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output110_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3279__I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output127_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output128_I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output137_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output146_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3294__I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output148_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3295__I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output162_I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output163_I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output164_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output165_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output166_I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output167_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3301__I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output168_I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output169_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output170_I (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3304__I (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output171_I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output174_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output175_I (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output186_I (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output187_I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output190_I (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output192_I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3306__I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output207_I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3310__I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output212_I (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output215_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3013__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3011__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3012__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__CLK (.I(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__CLK (.I(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__CLK (.I(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__CLK (.I(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2949__CLK (.I(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3147__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3143__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3043__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3133__CLK (.I(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2941__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3051__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3094__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3050__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2940__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3092__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3089__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3039__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2909__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3196__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__CLK (.I(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3076__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3041__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2914__CLK (.I(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3055__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3159__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3077__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3084__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3082__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3181__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3240__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3167__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__CLK (.I(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3063__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3245__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3244__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3243__CLK (.I(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3263__I (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__I (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3261__I (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3252__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__I (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3259__I (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3260__I (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3257__I (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3256__I (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3250__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3255__I (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3254__I (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3235__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2886__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3078__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3065__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3080__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__CLK (.I(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3074__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3069__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3072__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3073__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2972__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3079__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2975__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2907__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2977__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2979__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2922__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2851__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2982__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__CLK (.I(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2859__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2987__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2985__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2842__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2994__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2984__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2986__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2997__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3000__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2991__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3231__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3001__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2998__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2995__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3002__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3230__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2992__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2993__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3223__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2990__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2988__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2999__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2989__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2926__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3003__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3113__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3112__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3110__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3108__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3109__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3107__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3105__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3104__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2924__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3103__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3102__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3199__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3101__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2968__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2934__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3116__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3115__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3114__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3117__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3030__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3182__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3026__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3027__CLK (.I(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3025__CLK (.I(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3024__CLK (.I(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__CLK (.I(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2955__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2939__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3004__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2918__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3021__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3022__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3019__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3020__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3184__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3015__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3014__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3017__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3016__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3127__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3190__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_3__f_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_2__f_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_1__f_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_0__f_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_clock_I (.I(clknet_2_0__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_clock_I (.I(clknet_2_1__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_clock_I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_clock_I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_clock_I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_clock_I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_clock_I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_clock_I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_clock_I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_clock_I (.I(clknet_2_2__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_clock_I (.I(clknet_2_3__leaf_clock));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1399 ();
endmodule

