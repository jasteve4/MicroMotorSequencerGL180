// This is the unpowered netlist.
module driver_core (clock,
    clock_a,
    inverter_select_a,
    mem_write_n_a,
    output_active_a,
    row_col_select_a,
    col_select_a,
    data_in_a,
    driver_io,
    mem_address_a,
    row_select_a);
 input clock;
 input clock_a;
 input inverter_select_a;
 input mem_write_n_a;
 input output_active_a;
 input row_col_select_a;
 input [5:0] col_select_a;
 input [15:0] data_in_a;
 output [1:0] driver_io;
 input [9:0] mem_address_a;
 input [5:0] row_select_a;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire \col_select_trans[0].A ;
 wire \col_select_trans[0].data_sync ;
 wire \col_select_trans[1].A ;
 wire \col_select_trans[1].data_sync ;
 wire \col_select_trans[2].A ;
 wire \col_select_trans[2].data_sync ;
 wire \col_select_trans[3].A ;
 wire \col_select_trans[3].data_sync ;
 wire \col_select_trans[4].A ;
 wire \col_select_trans[4].data_sync ;
 wire \col_select_trans[5].A ;
 wire \col_select_trans[5].data_sync ;
 wire \data_in_trans[0].A ;
 wire \data_in_trans[0].data_sync ;
 wire \data_in_trans[10].A ;
 wire \data_in_trans[10].data_sync ;
 wire \data_in_trans[11].A ;
 wire \data_in_trans[11].data_sync ;
 wire \data_in_trans[12].A ;
 wire \data_in_trans[12].data_sync ;
 wire \data_in_trans[13].A ;
 wire \data_in_trans[13].data_sync ;
 wire \data_in_trans[14].A ;
 wire \data_in_trans[14].data_sync ;
 wire \data_in_trans[15].A ;
 wire \data_in_trans[15].data_sync ;
 wire \data_in_trans[1].A ;
 wire \data_in_trans[1].data_sync ;
 wire \data_in_trans[2].A ;
 wire \data_in_trans[2].data_sync ;
 wire \data_in_trans[3].A ;
 wire \data_in_trans[3].data_sync ;
 wire \data_in_trans[4].A ;
 wire \data_in_trans[4].data_sync ;
 wire \data_in_trans[5].A ;
 wire \data_in_trans[5].data_sync ;
 wire \data_in_trans[6].A ;
 wire \data_in_trans[6].data_sync ;
 wire \data_in_trans[7].A ;
 wire \data_in_trans[7].data_sync ;
 wire \data_in_trans[8].A ;
 wire \data_in_trans[8].data_sync ;
 wire \data_in_trans[9].A ;
 wire \data_in_trans[9].data_sync ;
 wire \inverter_select_trans.A ;
 wire \inverter_select_trans.data_sync ;
 wire \mem_address_trans[0].A ;
 wire \mem_address_trans[0].data_sync ;
 wire \mem_address_trans[1].A ;
 wire \mem_address_trans[1].data_sync ;
 wire \mem_address_trans[2].A ;
 wire \mem_address_trans[2].data_sync ;
 wire \mem_address_trans[3].A ;
 wire \mem_address_trans[3].data_sync ;
 wire \mem_address_trans[4].A ;
 wire \mem_address_trans[4].data_sync ;
 wire \mem_address_trans[5].A ;
 wire \mem_address_trans[5].data_sync ;
 wire \mem_address_trans[6].A ;
 wire \mem_address_trans[6].data_sync ;
 wire \mem_address_trans[7].A ;
 wire \mem_address_trans[7].data_sync ;
 wire \mem_address_trans[8].A ;
 wire \mem_address_trans[8].data_sync ;
 wire \mem_address_trans[9].A ;
 wire \mem_address_trans[9].data_sync ;
 wire \mem_write_n_trans.A ;
 wire \mem_write_n_trans.data_sync ;
 wire \output_active_hold[0] ;
 wire \output_active_hold[1] ;
 wire \output_active_hold[2] ;
 wire \output_active_hold[3] ;
 wire \output_active_trans.A ;
 wire \output_active_trans.data_sync ;
 wire \row_col_select_trans.A ;
 wire \row_col_select_trans.data_sync ;
 wire \row_select_trans[0].A ;
 wire \row_select_trans[0].data_sync ;
 wire \row_select_trans[1].A ;
 wire \row_select_trans[1].data_sync ;
 wire \row_select_trans[2].A ;
 wire \row_select_trans[2].data_sync ;
 wire \row_select_trans[3].A ;
 wire \row_select_trans[3].data_sync ;
 wire \row_select_trans[4].A ;
 wire \row_select_trans[4].data_sync ;
 wire \row_select_trans[5].A ;
 wire \row_select_trans[5].data_sync ;
 wire \u2.active_mem[0] ;
 wire \u2.active_mem[10] ;
 wire \u2.active_mem[11] ;
 wire \u2.active_mem[12] ;
 wire \u2.active_mem[13] ;
 wire \u2.active_mem[14] ;
 wire \u2.active_mem[15] ;
 wire \u2.active_mem[1] ;
 wire \u2.active_mem[2] ;
 wire \u2.active_mem[3] ;
 wire \u2.active_mem[4] ;
 wire \u2.active_mem[5] ;
 wire \u2.active_mem[6] ;
 wire \u2.active_mem[7] ;
 wire \u2.active_mem[8] ;
 wire \u2.active_mem[9] ;
 wire \u2.driver_enable ;
 wire \u2.driver_mem[0] ;
 wire \u2.driver_mem[10] ;
 wire \u2.driver_mem[11] ;
 wire \u2.driver_mem[12] ;
 wire \u2.driver_mem[13] ;
 wire \u2.driver_mem[14] ;
 wire \u2.driver_mem[15] ;
 wire \u2.driver_mem[1] ;
 wire \u2.driver_mem[2] ;
 wire \u2.driver_mem[3] ;
 wire \u2.driver_mem[4] ;
 wire \u2.driver_mem[5] ;
 wire \u2.driver_mem[6] ;
 wire \u2.driver_mem[7] ;
 wire \u2.driver_mem[8] ;
 wire \u2.driver_mem[9] ;
 wire \u2.mem[0][0] ;
 wire \u2.mem[0][10] ;
 wire \u2.mem[0][11] ;
 wire \u2.mem[0][12] ;
 wire \u2.mem[0][13] ;
 wire \u2.mem[0][14] ;
 wire \u2.mem[0][15] ;
 wire \u2.mem[0][1] ;
 wire \u2.mem[0][2] ;
 wire \u2.mem[0][3] ;
 wire \u2.mem[0][4] ;
 wire \u2.mem[0][5] ;
 wire \u2.mem[0][6] ;
 wire \u2.mem[0][7] ;
 wire \u2.mem[0][8] ;
 wire \u2.mem[0][9] ;
 wire \u2.mem[10][0] ;
 wire \u2.mem[10][10] ;
 wire \u2.mem[10][11] ;
 wire \u2.mem[10][12] ;
 wire \u2.mem[10][13] ;
 wire \u2.mem[10][14] ;
 wire \u2.mem[10][15] ;
 wire \u2.mem[10][1] ;
 wire \u2.mem[10][2] ;
 wire \u2.mem[10][3] ;
 wire \u2.mem[10][4] ;
 wire \u2.mem[10][5] ;
 wire \u2.mem[10][6] ;
 wire \u2.mem[10][7] ;
 wire \u2.mem[10][8] ;
 wire \u2.mem[10][9] ;
 wire \u2.mem[11][0] ;
 wire \u2.mem[11][10] ;
 wire \u2.mem[11][11] ;
 wire \u2.mem[11][12] ;
 wire \u2.mem[11][13] ;
 wire \u2.mem[11][14] ;
 wire \u2.mem[11][15] ;
 wire \u2.mem[11][1] ;
 wire \u2.mem[11][2] ;
 wire \u2.mem[11][3] ;
 wire \u2.mem[11][4] ;
 wire \u2.mem[11][5] ;
 wire \u2.mem[11][6] ;
 wire \u2.mem[11][7] ;
 wire \u2.mem[11][8] ;
 wire \u2.mem[11][9] ;
 wire \u2.mem[128][0] ;
 wire \u2.mem[128][1] ;
 wire \u2.mem[128][2] ;
 wire \u2.mem[128][3] ;
 wire \u2.mem[128][4] ;
 wire \u2.mem[128][5] ;
 wire \u2.mem[129][0] ;
 wire \u2.mem[129][1] ;
 wire \u2.mem[129][2] ;
 wire \u2.mem[129][3] ;
 wire \u2.mem[129][4] ;
 wire \u2.mem[129][5] ;
 wire \u2.mem[12][0] ;
 wire \u2.mem[12][10] ;
 wire \u2.mem[12][11] ;
 wire \u2.mem[12][12] ;
 wire \u2.mem[12][13] ;
 wire \u2.mem[12][14] ;
 wire \u2.mem[12][15] ;
 wire \u2.mem[12][1] ;
 wire \u2.mem[12][2] ;
 wire \u2.mem[12][3] ;
 wire \u2.mem[12][4] ;
 wire \u2.mem[12][5] ;
 wire \u2.mem[12][6] ;
 wire \u2.mem[12][7] ;
 wire \u2.mem[12][8] ;
 wire \u2.mem[12][9] ;
 wire \u2.mem[130][0] ;
 wire \u2.mem[130][1] ;
 wire \u2.mem[130][2] ;
 wire \u2.mem[130][3] ;
 wire \u2.mem[130][4] ;
 wire \u2.mem[130][5] ;
 wire \u2.mem[131][0] ;
 wire \u2.mem[131][1] ;
 wire \u2.mem[131][2] ;
 wire \u2.mem[131][3] ;
 wire \u2.mem[131][4] ;
 wire \u2.mem[131][5] ;
 wire \u2.mem[132][0] ;
 wire \u2.mem[132][1] ;
 wire \u2.mem[132][2] ;
 wire \u2.mem[132][3] ;
 wire \u2.mem[132][4] ;
 wire \u2.mem[132][5] ;
 wire \u2.mem[133][0] ;
 wire \u2.mem[133][1] ;
 wire \u2.mem[133][2] ;
 wire \u2.mem[133][3] ;
 wire \u2.mem[133][4] ;
 wire \u2.mem[133][5] ;
 wire \u2.mem[134][0] ;
 wire \u2.mem[134][1] ;
 wire \u2.mem[134][2] ;
 wire \u2.mem[134][3] ;
 wire \u2.mem[134][4] ;
 wire \u2.mem[134][5] ;
 wire \u2.mem[135][0] ;
 wire \u2.mem[135][1] ;
 wire \u2.mem[135][2] ;
 wire \u2.mem[135][3] ;
 wire \u2.mem[135][4] ;
 wire \u2.mem[135][5] ;
 wire \u2.mem[136][0] ;
 wire \u2.mem[136][1] ;
 wire \u2.mem[136][2] ;
 wire \u2.mem[136][3] ;
 wire \u2.mem[136][4] ;
 wire \u2.mem[136][5] ;
 wire \u2.mem[137][0] ;
 wire \u2.mem[137][1] ;
 wire \u2.mem[137][2] ;
 wire \u2.mem[137][3] ;
 wire \u2.mem[137][4] ;
 wire \u2.mem[137][5] ;
 wire \u2.mem[138][0] ;
 wire \u2.mem[138][1] ;
 wire \u2.mem[138][2] ;
 wire \u2.mem[138][3] ;
 wire \u2.mem[138][4] ;
 wire \u2.mem[138][5] ;
 wire \u2.mem[139][0] ;
 wire \u2.mem[139][1] ;
 wire \u2.mem[139][2] ;
 wire \u2.mem[139][3] ;
 wire \u2.mem[139][4] ;
 wire \u2.mem[139][5] ;
 wire \u2.mem[13][0] ;
 wire \u2.mem[13][10] ;
 wire \u2.mem[13][11] ;
 wire \u2.mem[13][12] ;
 wire \u2.mem[13][13] ;
 wire \u2.mem[13][14] ;
 wire \u2.mem[13][15] ;
 wire \u2.mem[13][1] ;
 wire \u2.mem[13][2] ;
 wire \u2.mem[13][3] ;
 wire \u2.mem[13][4] ;
 wire \u2.mem[13][5] ;
 wire \u2.mem[13][6] ;
 wire \u2.mem[13][7] ;
 wire \u2.mem[13][8] ;
 wire \u2.mem[13][9] ;
 wire \u2.mem[140][0] ;
 wire \u2.mem[140][1] ;
 wire \u2.mem[140][2] ;
 wire \u2.mem[140][3] ;
 wire \u2.mem[140][4] ;
 wire \u2.mem[140][5] ;
 wire \u2.mem[141][0] ;
 wire \u2.mem[141][1] ;
 wire \u2.mem[141][2] ;
 wire \u2.mem[141][3] ;
 wire \u2.mem[141][4] ;
 wire \u2.mem[141][5] ;
 wire \u2.mem[142][0] ;
 wire \u2.mem[142][1] ;
 wire \u2.mem[142][2] ;
 wire \u2.mem[142][3] ;
 wire \u2.mem[142][4] ;
 wire \u2.mem[142][5] ;
 wire \u2.mem[143][0] ;
 wire \u2.mem[143][1] ;
 wire \u2.mem[143][2] ;
 wire \u2.mem[143][3] ;
 wire \u2.mem[143][4] ;
 wire \u2.mem[143][5] ;
 wire \u2.mem[144][0] ;
 wire \u2.mem[144][1] ;
 wire \u2.mem[144][2] ;
 wire \u2.mem[144][3] ;
 wire \u2.mem[144][4] ;
 wire \u2.mem[144][5] ;
 wire \u2.mem[145][0] ;
 wire \u2.mem[145][1] ;
 wire \u2.mem[145][2] ;
 wire \u2.mem[145][3] ;
 wire \u2.mem[145][4] ;
 wire \u2.mem[145][5] ;
 wire \u2.mem[146][0] ;
 wire \u2.mem[146][1] ;
 wire \u2.mem[146][2] ;
 wire \u2.mem[146][3] ;
 wire \u2.mem[146][4] ;
 wire \u2.mem[146][5] ;
 wire \u2.mem[147][0] ;
 wire \u2.mem[147][1] ;
 wire \u2.mem[147][2] ;
 wire \u2.mem[147][3] ;
 wire \u2.mem[147][4] ;
 wire \u2.mem[147][5] ;
 wire \u2.mem[148][0] ;
 wire \u2.mem[148][1] ;
 wire \u2.mem[148][2] ;
 wire \u2.mem[148][3] ;
 wire \u2.mem[148][4] ;
 wire \u2.mem[148][5] ;
 wire \u2.mem[149][0] ;
 wire \u2.mem[149][1] ;
 wire \u2.mem[149][2] ;
 wire \u2.mem[149][3] ;
 wire \u2.mem[149][4] ;
 wire \u2.mem[149][5] ;
 wire \u2.mem[14][0] ;
 wire \u2.mem[14][10] ;
 wire \u2.mem[14][11] ;
 wire \u2.mem[14][12] ;
 wire \u2.mem[14][13] ;
 wire \u2.mem[14][14] ;
 wire \u2.mem[14][15] ;
 wire \u2.mem[14][1] ;
 wire \u2.mem[14][2] ;
 wire \u2.mem[14][3] ;
 wire \u2.mem[14][4] ;
 wire \u2.mem[14][5] ;
 wire \u2.mem[14][6] ;
 wire \u2.mem[14][7] ;
 wire \u2.mem[14][8] ;
 wire \u2.mem[14][9] ;
 wire \u2.mem[150][0] ;
 wire \u2.mem[150][1] ;
 wire \u2.mem[150][2] ;
 wire \u2.mem[150][3] ;
 wire \u2.mem[150][4] ;
 wire \u2.mem[150][5] ;
 wire \u2.mem[151][0] ;
 wire \u2.mem[151][1] ;
 wire \u2.mem[151][2] ;
 wire \u2.mem[151][3] ;
 wire \u2.mem[151][4] ;
 wire \u2.mem[151][5] ;
 wire \u2.mem[152][0] ;
 wire \u2.mem[152][1] ;
 wire \u2.mem[152][2] ;
 wire \u2.mem[152][3] ;
 wire \u2.mem[152][4] ;
 wire \u2.mem[152][5] ;
 wire \u2.mem[153][0] ;
 wire \u2.mem[153][1] ;
 wire \u2.mem[153][2] ;
 wire \u2.mem[153][3] ;
 wire \u2.mem[153][4] ;
 wire \u2.mem[153][5] ;
 wire \u2.mem[154][0] ;
 wire \u2.mem[154][1] ;
 wire \u2.mem[154][2] ;
 wire \u2.mem[154][3] ;
 wire \u2.mem[154][4] ;
 wire \u2.mem[154][5] ;
 wire \u2.mem[155][0] ;
 wire \u2.mem[155][1] ;
 wire \u2.mem[155][2] ;
 wire \u2.mem[155][3] ;
 wire \u2.mem[155][4] ;
 wire \u2.mem[155][5] ;
 wire \u2.mem[156][0] ;
 wire \u2.mem[156][1] ;
 wire \u2.mem[156][2] ;
 wire \u2.mem[156][3] ;
 wire \u2.mem[156][4] ;
 wire \u2.mem[156][5] ;
 wire \u2.mem[157][0] ;
 wire \u2.mem[157][1] ;
 wire \u2.mem[157][2] ;
 wire \u2.mem[157][3] ;
 wire \u2.mem[157][4] ;
 wire \u2.mem[157][5] ;
 wire \u2.mem[158][0] ;
 wire \u2.mem[158][1] ;
 wire \u2.mem[158][2] ;
 wire \u2.mem[158][3] ;
 wire \u2.mem[158][4] ;
 wire \u2.mem[158][5] ;
 wire \u2.mem[159][0] ;
 wire \u2.mem[159][1] ;
 wire \u2.mem[159][2] ;
 wire \u2.mem[159][3] ;
 wire \u2.mem[159][4] ;
 wire \u2.mem[159][5] ;
 wire \u2.mem[15][0] ;
 wire \u2.mem[15][10] ;
 wire \u2.mem[15][11] ;
 wire \u2.mem[15][12] ;
 wire \u2.mem[15][13] ;
 wire \u2.mem[15][14] ;
 wire \u2.mem[15][15] ;
 wire \u2.mem[15][1] ;
 wire \u2.mem[15][2] ;
 wire \u2.mem[15][3] ;
 wire \u2.mem[15][4] ;
 wire \u2.mem[15][5] ;
 wire \u2.mem[15][6] ;
 wire \u2.mem[15][7] ;
 wire \u2.mem[15][8] ;
 wire \u2.mem[15][9] ;
 wire \u2.mem[160][0] ;
 wire \u2.mem[160][1] ;
 wire \u2.mem[160][2] ;
 wire \u2.mem[160][3] ;
 wire \u2.mem[160][4] ;
 wire \u2.mem[160][5] ;
 wire \u2.mem[161][0] ;
 wire \u2.mem[161][1] ;
 wire \u2.mem[161][2] ;
 wire \u2.mem[161][3] ;
 wire \u2.mem[161][4] ;
 wire \u2.mem[161][5] ;
 wire \u2.mem[162][0] ;
 wire \u2.mem[162][1] ;
 wire \u2.mem[162][2] ;
 wire \u2.mem[162][3] ;
 wire \u2.mem[162][4] ;
 wire \u2.mem[162][5] ;
 wire \u2.mem[163][0] ;
 wire \u2.mem[163][1] ;
 wire \u2.mem[163][2] ;
 wire \u2.mem[163][3] ;
 wire \u2.mem[163][4] ;
 wire \u2.mem[163][5] ;
 wire \u2.mem[164][0] ;
 wire \u2.mem[164][1] ;
 wire \u2.mem[164][2] ;
 wire \u2.mem[164][3] ;
 wire \u2.mem[164][4] ;
 wire \u2.mem[164][5] ;
 wire \u2.mem[165][0] ;
 wire \u2.mem[165][1] ;
 wire \u2.mem[165][2] ;
 wire \u2.mem[165][3] ;
 wire \u2.mem[165][4] ;
 wire \u2.mem[165][5] ;
 wire \u2.mem[166][0] ;
 wire \u2.mem[166][1] ;
 wire \u2.mem[166][2] ;
 wire \u2.mem[166][3] ;
 wire \u2.mem[166][4] ;
 wire \u2.mem[166][5] ;
 wire \u2.mem[167][0] ;
 wire \u2.mem[167][1] ;
 wire \u2.mem[167][2] ;
 wire \u2.mem[167][3] ;
 wire \u2.mem[167][4] ;
 wire \u2.mem[167][5] ;
 wire \u2.mem[168][0] ;
 wire \u2.mem[168][1] ;
 wire \u2.mem[168][2] ;
 wire \u2.mem[168][3] ;
 wire \u2.mem[168][4] ;
 wire \u2.mem[168][5] ;
 wire \u2.mem[169][0] ;
 wire \u2.mem[169][1] ;
 wire \u2.mem[169][2] ;
 wire \u2.mem[169][3] ;
 wire \u2.mem[169][4] ;
 wire \u2.mem[169][5] ;
 wire \u2.mem[16][0] ;
 wire \u2.mem[16][10] ;
 wire \u2.mem[16][11] ;
 wire \u2.mem[16][12] ;
 wire \u2.mem[16][13] ;
 wire \u2.mem[16][14] ;
 wire \u2.mem[16][15] ;
 wire \u2.mem[16][1] ;
 wire \u2.mem[16][2] ;
 wire \u2.mem[16][3] ;
 wire \u2.mem[16][4] ;
 wire \u2.mem[16][5] ;
 wire \u2.mem[16][6] ;
 wire \u2.mem[16][7] ;
 wire \u2.mem[16][8] ;
 wire \u2.mem[16][9] ;
 wire \u2.mem[170][0] ;
 wire \u2.mem[170][1] ;
 wire \u2.mem[170][2] ;
 wire \u2.mem[170][3] ;
 wire \u2.mem[170][4] ;
 wire \u2.mem[170][5] ;
 wire \u2.mem[171][0] ;
 wire \u2.mem[171][1] ;
 wire \u2.mem[171][2] ;
 wire \u2.mem[171][3] ;
 wire \u2.mem[171][4] ;
 wire \u2.mem[171][5] ;
 wire \u2.mem[172][0] ;
 wire \u2.mem[172][1] ;
 wire \u2.mem[172][2] ;
 wire \u2.mem[172][3] ;
 wire \u2.mem[172][4] ;
 wire \u2.mem[172][5] ;
 wire \u2.mem[173][0] ;
 wire \u2.mem[173][1] ;
 wire \u2.mem[173][2] ;
 wire \u2.mem[173][3] ;
 wire \u2.mem[173][4] ;
 wire \u2.mem[173][5] ;
 wire \u2.mem[174][0] ;
 wire \u2.mem[174][1] ;
 wire \u2.mem[174][2] ;
 wire \u2.mem[174][3] ;
 wire \u2.mem[174][4] ;
 wire \u2.mem[174][5] ;
 wire \u2.mem[175][0] ;
 wire \u2.mem[175][1] ;
 wire \u2.mem[175][2] ;
 wire \u2.mem[175][3] ;
 wire \u2.mem[175][4] ;
 wire \u2.mem[175][5] ;
 wire \u2.mem[176][0] ;
 wire \u2.mem[176][1] ;
 wire \u2.mem[176][2] ;
 wire \u2.mem[176][3] ;
 wire \u2.mem[176][4] ;
 wire \u2.mem[176][5] ;
 wire \u2.mem[177][0] ;
 wire \u2.mem[177][1] ;
 wire \u2.mem[177][2] ;
 wire \u2.mem[177][3] ;
 wire \u2.mem[177][4] ;
 wire \u2.mem[177][5] ;
 wire \u2.mem[178][0] ;
 wire \u2.mem[178][1] ;
 wire \u2.mem[178][2] ;
 wire \u2.mem[178][3] ;
 wire \u2.mem[178][4] ;
 wire \u2.mem[178][5] ;
 wire \u2.mem[179][0] ;
 wire \u2.mem[179][1] ;
 wire \u2.mem[179][2] ;
 wire \u2.mem[179][3] ;
 wire \u2.mem[179][4] ;
 wire \u2.mem[179][5] ;
 wire \u2.mem[17][0] ;
 wire \u2.mem[17][10] ;
 wire \u2.mem[17][11] ;
 wire \u2.mem[17][12] ;
 wire \u2.mem[17][13] ;
 wire \u2.mem[17][14] ;
 wire \u2.mem[17][15] ;
 wire \u2.mem[17][1] ;
 wire \u2.mem[17][2] ;
 wire \u2.mem[17][3] ;
 wire \u2.mem[17][4] ;
 wire \u2.mem[17][5] ;
 wire \u2.mem[17][6] ;
 wire \u2.mem[17][7] ;
 wire \u2.mem[17][8] ;
 wire \u2.mem[17][9] ;
 wire \u2.mem[180][0] ;
 wire \u2.mem[180][1] ;
 wire \u2.mem[180][2] ;
 wire \u2.mem[180][3] ;
 wire \u2.mem[180][4] ;
 wire \u2.mem[180][5] ;
 wire \u2.mem[181][0] ;
 wire \u2.mem[181][1] ;
 wire \u2.mem[181][2] ;
 wire \u2.mem[181][3] ;
 wire \u2.mem[181][4] ;
 wire \u2.mem[181][5] ;
 wire \u2.mem[182][0] ;
 wire \u2.mem[182][1] ;
 wire \u2.mem[182][2] ;
 wire \u2.mem[182][3] ;
 wire \u2.mem[182][4] ;
 wire \u2.mem[182][5] ;
 wire \u2.mem[183][0] ;
 wire \u2.mem[183][1] ;
 wire \u2.mem[183][2] ;
 wire \u2.mem[183][3] ;
 wire \u2.mem[183][4] ;
 wire \u2.mem[183][5] ;
 wire \u2.mem[184][0] ;
 wire \u2.mem[184][1] ;
 wire \u2.mem[184][2] ;
 wire \u2.mem[184][3] ;
 wire \u2.mem[184][4] ;
 wire \u2.mem[184][5] ;
 wire \u2.mem[185][0] ;
 wire \u2.mem[185][1] ;
 wire \u2.mem[185][2] ;
 wire \u2.mem[185][3] ;
 wire \u2.mem[185][4] ;
 wire \u2.mem[185][5] ;
 wire \u2.mem[186][0] ;
 wire \u2.mem[186][1] ;
 wire \u2.mem[186][2] ;
 wire \u2.mem[186][3] ;
 wire \u2.mem[186][4] ;
 wire \u2.mem[186][5] ;
 wire \u2.mem[187][0] ;
 wire \u2.mem[187][1] ;
 wire \u2.mem[187][2] ;
 wire \u2.mem[187][3] ;
 wire \u2.mem[187][4] ;
 wire \u2.mem[187][5] ;
 wire \u2.mem[188][0] ;
 wire \u2.mem[188][1] ;
 wire \u2.mem[188][2] ;
 wire \u2.mem[188][3] ;
 wire \u2.mem[188][4] ;
 wire \u2.mem[188][5] ;
 wire \u2.mem[189][0] ;
 wire \u2.mem[189][1] ;
 wire \u2.mem[189][2] ;
 wire \u2.mem[189][3] ;
 wire \u2.mem[189][4] ;
 wire \u2.mem[189][5] ;
 wire \u2.mem[18][0] ;
 wire \u2.mem[18][10] ;
 wire \u2.mem[18][11] ;
 wire \u2.mem[18][12] ;
 wire \u2.mem[18][13] ;
 wire \u2.mem[18][14] ;
 wire \u2.mem[18][15] ;
 wire \u2.mem[18][1] ;
 wire \u2.mem[18][2] ;
 wire \u2.mem[18][3] ;
 wire \u2.mem[18][4] ;
 wire \u2.mem[18][5] ;
 wire \u2.mem[18][6] ;
 wire \u2.mem[18][7] ;
 wire \u2.mem[18][8] ;
 wire \u2.mem[18][9] ;
 wire \u2.mem[190][0] ;
 wire \u2.mem[190][1] ;
 wire \u2.mem[190][2] ;
 wire \u2.mem[190][3] ;
 wire \u2.mem[190][4] ;
 wire \u2.mem[190][5] ;
 wire \u2.mem[191][0] ;
 wire \u2.mem[191][1] ;
 wire \u2.mem[191][2] ;
 wire \u2.mem[191][3] ;
 wire \u2.mem[191][4] ;
 wire \u2.mem[191][5] ;
 wire \u2.mem[192][0] ;
 wire \u2.mem[192][10] ;
 wire \u2.mem[192][11] ;
 wire \u2.mem[192][12] ;
 wire \u2.mem[192][13] ;
 wire \u2.mem[192][14] ;
 wire \u2.mem[192][15] ;
 wire \u2.mem[192][1] ;
 wire \u2.mem[192][2] ;
 wire \u2.mem[192][3] ;
 wire \u2.mem[192][4] ;
 wire \u2.mem[192][5] ;
 wire \u2.mem[192][6] ;
 wire \u2.mem[192][7] ;
 wire \u2.mem[192][8] ;
 wire \u2.mem[192][9] ;
 wire \u2.mem[193][0] ;
 wire \u2.mem[193][10] ;
 wire \u2.mem[193][11] ;
 wire \u2.mem[193][12] ;
 wire \u2.mem[193][13] ;
 wire \u2.mem[193][14] ;
 wire \u2.mem[193][15] ;
 wire \u2.mem[193][1] ;
 wire \u2.mem[193][2] ;
 wire \u2.mem[193][3] ;
 wire \u2.mem[193][4] ;
 wire \u2.mem[193][5] ;
 wire \u2.mem[193][6] ;
 wire \u2.mem[193][7] ;
 wire \u2.mem[193][8] ;
 wire \u2.mem[193][9] ;
 wire \u2.mem[194][0] ;
 wire \u2.mem[194][10] ;
 wire \u2.mem[194][11] ;
 wire \u2.mem[194][12] ;
 wire \u2.mem[194][13] ;
 wire \u2.mem[194][14] ;
 wire \u2.mem[194][15] ;
 wire \u2.mem[194][1] ;
 wire \u2.mem[194][2] ;
 wire \u2.mem[194][3] ;
 wire \u2.mem[194][4] ;
 wire \u2.mem[194][5] ;
 wire \u2.mem[194][6] ;
 wire \u2.mem[194][7] ;
 wire \u2.mem[194][8] ;
 wire \u2.mem[194][9] ;
 wire \u2.mem[19][0] ;
 wire \u2.mem[19][10] ;
 wire \u2.mem[19][11] ;
 wire \u2.mem[19][12] ;
 wire \u2.mem[19][13] ;
 wire \u2.mem[19][14] ;
 wire \u2.mem[19][15] ;
 wire \u2.mem[19][1] ;
 wire \u2.mem[19][2] ;
 wire \u2.mem[19][3] ;
 wire \u2.mem[19][4] ;
 wire \u2.mem[19][5] ;
 wire \u2.mem[19][6] ;
 wire \u2.mem[19][7] ;
 wire \u2.mem[19][8] ;
 wire \u2.mem[19][9] ;
 wire \u2.mem[1][0] ;
 wire \u2.mem[1][10] ;
 wire \u2.mem[1][11] ;
 wire \u2.mem[1][12] ;
 wire \u2.mem[1][13] ;
 wire \u2.mem[1][14] ;
 wire \u2.mem[1][15] ;
 wire \u2.mem[1][1] ;
 wire \u2.mem[1][2] ;
 wire \u2.mem[1][3] ;
 wire \u2.mem[1][4] ;
 wire \u2.mem[1][5] ;
 wire \u2.mem[1][6] ;
 wire \u2.mem[1][7] ;
 wire \u2.mem[1][8] ;
 wire \u2.mem[1][9] ;
 wire \u2.mem[20][0] ;
 wire \u2.mem[20][10] ;
 wire \u2.mem[20][11] ;
 wire \u2.mem[20][12] ;
 wire \u2.mem[20][13] ;
 wire \u2.mem[20][14] ;
 wire \u2.mem[20][15] ;
 wire \u2.mem[20][1] ;
 wire \u2.mem[20][2] ;
 wire \u2.mem[20][3] ;
 wire \u2.mem[20][4] ;
 wire \u2.mem[20][5] ;
 wire \u2.mem[20][6] ;
 wire \u2.mem[20][7] ;
 wire \u2.mem[20][8] ;
 wire \u2.mem[20][9] ;
 wire \u2.mem[21][0] ;
 wire \u2.mem[21][10] ;
 wire \u2.mem[21][11] ;
 wire \u2.mem[21][12] ;
 wire \u2.mem[21][13] ;
 wire \u2.mem[21][14] ;
 wire \u2.mem[21][15] ;
 wire \u2.mem[21][1] ;
 wire \u2.mem[21][2] ;
 wire \u2.mem[21][3] ;
 wire \u2.mem[21][4] ;
 wire \u2.mem[21][5] ;
 wire \u2.mem[21][6] ;
 wire \u2.mem[21][7] ;
 wire \u2.mem[21][8] ;
 wire \u2.mem[21][9] ;
 wire \u2.mem[22][0] ;
 wire \u2.mem[22][10] ;
 wire \u2.mem[22][11] ;
 wire \u2.mem[22][12] ;
 wire \u2.mem[22][13] ;
 wire \u2.mem[22][14] ;
 wire \u2.mem[22][15] ;
 wire \u2.mem[22][1] ;
 wire \u2.mem[22][2] ;
 wire \u2.mem[22][3] ;
 wire \u2.mem[22][4] ;
 wire \u2.mem[22][5] ;
 wire \u2.mem[22][6] ;
 wire \u2.mem[22][7] ;
 wire \u2.mem[22][8] ;
 wire \u2.mem[22][9] ;
 wire \u2.mem[23][0] ;
 wire \u2.mem[23][10] ;
 wire \u2.mem[23][11] ;
 wire \u2.mem[23][12] ;
 wire \u2.mem[23][13] ;
 wire \u2.mem[23][14] ;
 wire \u2.mem[23][15] ;
 wire \u2.mem[23][1] ;
 wire \u2.mem[23][2] ;
 wire \u2.mem[23][3] ;
 wire \u2.mem[23][4] ;
 wire \u2.mem[23][5] ;
 wire \u2.mem[23][6] ;
 wire \u2.mem[23][7] ;
 wire \u2.mem[23][8] ;
 wire \u2.mem[23][9] ;
 wire \u2.mem[24][0] ;
 wire \u2.mem[24][10] ;
 wire \u2.mem[24][11] ;
 wire \u2.mem[24][12] ;
 wire \u2.mem[24][13] ;
 wire \u2.mem[24][14] ;
 wire \u2.mem[24][15] ;
 wire \u2.mem[24][1] ;
 wire \u2.mem[24][2] ;
 wire \u2.mem[24][3] ;
 wire \u2.mem[24][4] ;
 wire \u2.mem[24][5] ;
 wire \u2.mem[24][6] ;
 wire \u2.mem[24][7] ;
 wire \u2.mem[24][8] ;
 wire \u2.mem[24][9] ;
 wire \u2.mem[25][0] ;
 wire \u2.mem[25][10] ;
 wire \u2.mem[25][11] ;
 wire \u2.mem[25][12] ;
 wire \u2.mem[25][13] ;
 wire \u2.mem[25][14] ;
 wire \u2.mem[25][15] ;
 wire \u2.mem[25][1] ;
 wire \u2.mem[25][2] ;
 wire \u2.mem[25][3] ;
 wire \u2.mem[25][4] ;
 wire \u2.mem[25][5] ;
 wire \u2.mem[25][6] ;
 wire \u2.mem[25][7] ;
 wire \u2.mem[25][8] ;
 wire \u2.mem[25][9] ;
 wire \u2.mem[26][0] ;
 wire \u2.mem[26][10] ;
 wire \u2.mem[26][11] ;
 wire \u2.mem[26][12] ;
 wire \u2.mem[26][13] ;
 wire \u2.mem[26][14] ;
 wire \u2.mem[26][15] ;
 wire \u2.mem[26][1] ;
 wire \u2.mem[26][2] ;
 wire \u2.mem[26][3] ;
 wire \u2.mem[26][4] ;
 wire \u2.mem[26][5] ;
 wire \u2.mem[26][6] ;
 wire \u2.mem[26][7] ;
 wire \u2.mem[26][8] ;
 wire \u2.mem[26][9] ;
 wire \u2.mem[27][0] ;
 wire \u2.mem[27][10] ;
 wire \u2.mem[27][11] ;
 wire \u2.mem[27][12] ;
 wire \u2.mem[27][13] ;
 wire \u2.mem[27][14] ;
 wire \u2.mem[27][15] ;
 wire \u2.mem[27][1] ;
 wire \u2.mem[27][2] ;
 wire \u2.mem[27][3] ;
 wire \u2.mem[27][4] ;
 wire \u2.mem[27][5] ;
 wire \u2.mem[27][6] ;
 wire \u2.mem[27][7] ;
 wire \u2.mem[27][8] ;
 wire \u2.mem[27][9] ;
 wire \u2.mem[28][0] ;
 wire \u2.mem[28][10] ;
 wire \u2.mem[28][11] ;
 wire \u2.mem[28][12] ;
 wire \u2.mem[28][13] ;
 wire \u2.mem[28][14] ;
 wire \u2.mem[28][15] ;
 wire \u2.mem[28][1] ;
 wire \u2.mem[28][2] ;
 wire \u2.mem[28][3] ;
 wire \u2.mem[28][4] ;
 wire \u2.mem[28][5] ;
 wire \u2.mem[28][6] ;
 wire \u2.mem[28][7] ;
 wire \u2.mem[28][8] ;
 wire \u2.mem[28][9] ;
 wire \u2.mem[29][0] ;
 wire \u2.mem[29][10] ;
 wire \u2.mem[29][11] ;
 wire \u2.mem[29][12] ;
 wire \u2.mem[29][13] ;
 wire \u2.mem[29][14] ;
 wire \u2.mem[29][15] ;
 wire \u2.mem[29][1] ;
 wire \u2.mem[29][2] ;
 wire \u2.mem[29][3] ;
 wire \u2.mem[29][4] ;
 wire \u2.mem[29][5] ;
 wire \u2.mem[29][6] ;
 wire \u2.mem[29][7] ;
 wire \u2.mem[29][8] ;
 wire \u2.mem[29][9] ;
 wire \u2.mem[2][0] ;
 wire \u2.mem[2][10] ;
 wire \u2.mem[2][11] ;
 wire \u2.mem[2][12] ;
 wire \u2.mem[2][13] ;
 wire \u2.mem[2][14] ;
 wire \u2.mem[2][15] ;
 wire \u2.mem[2][1] ;
 wire \u2.mem[2][2] ;
 wire \u2.mem[2][3] ;
 wire \u2.mem[2][4] ;
 wire \u2.mem[2][5] ;
 wire \u2.mem[2][6] ;
 wire \u2.mem[2][7] ;
 wire \u2.mem[2][8] ;
 wire \u2.mem[2][9] ;
 wire \u2.mem[30][0] ;
 wire \u2.mem[30][10] ;
 wire \u2.mem[30][11] ;
 wire \u2.mem[30][12] ;
 wire \u2.mem[30][13] ;
 wire \u2.mem[30][14] ;
 wire \u2.mem[30][15] ;
 wire \u2.mem[30][1] ;
 wire \u2.mem[30][2] ;
 wire \u2.mem[30][3] ;
 wire \u2.mem[30][4] ;
 wire \u2.mem[30][5] ;
 wire \u2.mem[30][6] ;
 wire \u2.mem[30][7] ;
 wire \u2.mem[30][8] ;
 wire \u2.mem[30][9] ;
 wire \u2.mem[31][0] ;
 wire \u2.mem[31][10] ;
 wire \u2.mem[31][11] ;
 wire \u2.mem[31][12] ;
 wire \u2.mem[31][13] ;
 wire \u2.mem[31][14] ;
 wire \u2.mem[31][15] ;
 wire \u2.mem[31][1] ;
 wire \u2.mem[31][2] ;
 wire \u2.mem[31][3] ;
 wire \u2.mem[31][4] ;
 wire \u2.mem[31][5] ;
 wire \u2.mem[31][6] ;
 wire \u2.mem[31][7] ;
 wire \u2.mem[31][8] ;
 wire \u2.mem[31][9] ;
 wire \u2.mem[32][0] ;
 wire \u2.mem[32][10] ;
 wire \u2.mem[32][11] ;
 wire \u2.mem[32][12] ;
 wire \u2.mem[32][13] ;
 wire \u2.mem[32][14] ;
 wire \u2.mem[32][15] ;
 wire \u2.mem[32][1] ;
 wire \u2.mem[32][2] ;
 wire \u2.mem[32][3] ;
 wire \u2.mem[32][4] ;
 wire \u2.mem[32][5] ;
 wire \u2.mem[32][6] ;
 wire \u2.mem[32][7] ;
 wire \u2.mem[32][8] ;
 wire \u2.mem[32][9] ;
 wire \u2.mem[33][0] ;
 wire \u2.mem[33][10] ;
 wire \u2.mem[33][11] ;
 wire \u2.mem[33][12] ;
 wire \u2.mem[33][13] ;
 wire \u2.mem[33][14] ;
 wire \u2.mem[33][15] ;
 wire \u2.mem[33][1] ;
 wire \u2.mem[33][2] ;
 wire \u2.mem[33][3] ;
 wire \u2.mem[33][4] ;
 wire \u2.mem[33][5] ;
 wire \u2.mem[33][6] ;
 wire \u2.mem[33][7] ;
 wire \u2.mem[33][8] ;
 wire \u2.mem[33][9] ;
 wire \u2.mem[34][0] ;
 wire \u2.mem[34][10] ;
 wire \u2.mem[34][11] ;
 wire \u2.mem[34][12] ;
 wire \u2.mem[34][13] ;
 wire \u2.mem[34][14] ;
 wire \u2.mem[34][15] ;
 wire \u2.mem[34][1] ;
 wire \u2.mem[34][2] ;
 wire \u2.mem[34][3] ;
 wire \u2.mem[34][4] ;
 wire \u2.mem[34][5] ;
 wire \u2.mem[34][6] ;
 wire \u2.mem[34][7] ;
 wire \u2.mem[34][8] ;
 wire \u2.mem[34][9] ;
 wire \u2.mem[35][0] ;
 wire \u2.mem[35][10] ;
 wire \u2.mem[35][11] ;
 wire \u2.mem[35][12] ;
 wire \u2.mem[35][13] ;
 wire \u2.mem[35][14] ;
 wire \u2.mem[35][15] ;
 wire \u2.mem[35][1] ;
 wire \u2.mem[35][2] ;
 wire \u2.mem[35][3] ;
 wire \u2.mem[35][4] ;
 wire \u2.mem[35][5] ;
 wire \u2.mem[35][6] ;
 wire \u2.mem[35][7] ;
 wire \u2.mem[35][8] ;
 wire \u2.mem[35][9] ;
 wire \u2.mem[36][0] ;
 wire \u2.mem[36][10] ;
 wire \u2.mem[36][11] ;
 wire \u2.mem[36][12] ;
 wire \u2.mem[36][13] ;
 wire \u2.mem[36][14] ;
 wire \u2.mem[36][15] ;
 wire \u2.mem[36][1] ;
 wire \u2.mem[36][2] ;
 wire \u2.mem[36][3] ;
 wire \u2.mem[36][4] ;
 wire \u2.mem[36][5] ;
 wire \u2.mem[36][6] ;
 wire \u2.mem[36][7] ;
 wire \u2.mem[36][8] ;
 wire \u2.mem[36][9] ;
 wire \u2.mem[37][0] ;
 wire \u2.mem[37][10] ;
 wire \u2.mem[37][11] ;
 wire \u2.mem[37][12] ;
 wire \u2.mem[37][13] ;
 wire \u2.mem[37][14] ;
 wire \u2.mem[37][15] ;
 wire \u2.mem[37][1] ;
 wire \u2.mem[37][2] ;
 wire \u2.mem[37][3] ;
 wire \u2.mem[37][4] ;
 wire \u2.mem[37][5] ;
 wire \u2.mem[37][6] ;
 wire \u2.mem[37][7] ;
 wire \u2.mem[37][8] ;
 wire \u2.mem[37][9] ;
 wire \u2.mem[38][0] ;
 wire \u2.mem[38][10] ;
 wire \u2.mem[38][11] ;
 wire \u2.mem[38][12] ;
 wire \u2.mem[38][13] ;
 wire \u2.mem[38][14] ;
 wire \u2.mem[38][15] ;
 wire \u2.mem[38][1] ;
 wire \u2.mem[38][2] ;
 wire \u2.mem[38][3] ;
 wire \u2.mem[38][4] ;
 wire \u2.mem[38][5] ;
 wire \u2.mem[38][6] ;
 wire \u2.mem[38][7] ;
 wire \u2.mem[38][8] ;
 wire \u2.mem[38][9] ;
 wire \u2.mem[39][0] ;
 wire \u2.mem[39][10] ;
 wire \u2.mem[39][11] ;
 wire \u2.mem[39][12] ;
 wire \u2.mem[39][13] ;
 wire \u2.mem[39][14] ;
 wire \u2.mem[39][15] ;
 wire \u2.mem[39][1] ;
 wire \u2.mem[39][2] ;
 wire \u2.mem[39][3] ;
 wire \u2.mem[39][4] ;
 wire \u2.mem[39][5] ;
 wire \u2.mem[39][6] ;
 wire \u2.mem[39][7] ;
 wire \u2.mem[39][8] ;
 wire \u2.mem[39][9] ;
 wire \u2.mem[3][0] ;
 wire \u2.mem[3][10] ;
 wire \u2.mem[3][11] ;
 wire \u2.mem[3][12] ;
 wire \u2.mem[3][13] ;
 wire \u2.mem[3][14] ;
 wire \u2.mem[3][15] ;
 wire \u2.mem[3][1] ;
 wire \u2.mem[3][2] ;
 wire \u2.mem[3][3] ;
 wire \u2.mem[3][4] ;
 wire \u2.mem[3][5] ;
 wire \u2.mem[3][6] ;
 wire \u2.mem[3][7] ;
 wire \u2.mem[3][8] ;
 wire \u2.mem[3][9] ;
 wire \u2.mem[40][0] ;
 wire \u2.mem[40][10] ;
 wire \u2.mem[40][11] ;
 wire \u2.mem[40][12] ;
 wire \u2.mem[40][13] ;
 wire \u2.mem[40][14] ;
 wire \u2.mem[40][15] ;
 wire \u2.mem[40][1] ;
 wire \u2.mem[40][2] ;
 wire \u2.mem[40][3] ;
 wire \u2.mem[40][4] ;
 wire \u2.mem[40][5] ;
 wire \u2.mem[40][6] ;
 wire \u2.mem[40][7] ;
 wire \u2.mem[40][8] ;
 wire \u2.mem[40][9] ;
 wire \u2.mem[41][0] ;
 wire \u2.mem[41][10] ;
 wire \u2.mem[41][11] ;
 wire \u2.mem[41][12] ;
 wire \u2.mem[41][13] ;
 wire \u2.mem[41][14] ;
 wire \u2.mem[41][15] ;
 wire \u2.mem[41][1] ;
 wire \u2.mem[41][2] ;
 wire \u2.mem[41][3] ;
 wire \u2.mem[41][4] ;
 wire \u2.mem[41][5] ;
 wire \u2.mem[41][6] ;
 wire \u2.mem[41][7] ;
 wire \u2.mem[41][8] ;
 wire \u2.mem[41][9] ;
 wire \u2.mem[42][0] ;
 wire \u2.mem[42][10] ;
 wire \u2.mem[42][11] ;
 wire \u2.mem[42][12] ;
 wire \u2.mem[42][13] ;
 wire \u2.mem[42][14] ;
 wire \u2.mem[42][15] ;
 wire \u2.mem[42][1] ;
 wire \u2.mem[42][2] ;
 wire \u2.mem[42][3] ;
 wire \u2.mem[42][4] ;
 wire \u2.mem[42][5] ;
 wire \u2.mem[42][6] ;
 wire \u2.mem[42][7] ;
 wire \u2.mem[42][8] ;
 wire \u2.mem[42][9] ;
 wire \u2.mem[43][0] ;
 wire \u2.mem[43][10] ;
 wire \u2.mem[43][11] ;
 wire \u2.mem[43][12] ;
 wire \u2.mem[43][13] ;
 wire \u2.mem[43][14] ;
 wire \u2.mem[43][15] ;
 wire \u2.mem[43][1] ;
 wire \u2.mem[43][2] ;
 wire \u2.mem[43][3] ;
 wire \u2.mem[43][4] ;
 wire \u2.mem[43][5] ;
 wire \u2.mem[43][6] ;
 wire \u2.mem[43][7] ;
 wire \u2.mem[43][8] ;
 wire \u2.mem[43][9] ;
 wire \u2.mem[44][0] ;
 wire \u2.mem[44][10] ;
 wire \u2.mem[44][11] ;
 wire \u2.mem[44][12] ;
 wire \u2.mem[44][13] ;
 wire \u2.mem[44][14] ;
 wire \u2.mem[44][15] ;
 wire \u2.mem[44][1] ;
 wire \u2.mem[44][2] ;
 wire \u2.mem[44][3] ;
 wire \u2.mem[44][4] ;
 wire \u2.mem[44][5] ;
 wire \u2.mem[44][6] ;
 wire \u2.mem[44][7] ;
 wire \u2.mem[44][8] ;
 wire \u2.mem[44][9] ;
 wire \u2.mem[45][0] ;
 wire \u2.mem[45][10] ;
 wire \u2.mem[45][11] ;
 wire \u2.mem[45][12] ;
 wire \u2.mem[45][13] ;
 wire \u2.mem[45][14] ;
 wire \u2.mem[45][15] ;
 wire \u2.mem[45][1] ;
 wire \u2.mem[45][2] ;
 wire \u2.mem[45][3] ;
 wire \u2.mem[45][4] ;
 wire \u2.mem[45][5] ;
 wire \u2.mem[45][6] ;
 wire \u2.mem[45][7] ;
 wire \u2.mem[45][8] ;
 wire \u2.mem[45][9] ;
 wire \u2.mem[46][0] ;
 wire \u2.mem[46][10] ;
 wire \u2.mem[46][11] ;
 wire \u2.mem[46][12] ;
 wire \u2.mem[46][13] ;
 wire \u2.mem[46][14] ;
 wire \u2.mem[46][15] ;
 wire \u2.mem[46][1] ;
 wire \u2.mem[46][2] ;
 wire \u2.mem[46][3] ;
 wire \u2.mem[46][4] ;
 wire \u2.mem[46][5] ;
 wire \u2.mem[46][6] ;
 wire \u2.mem[46][7] ;
 wire \u2.mem[46][8] ;
 wire \u2.mem[46][9] ;
 wire \u2.mem[47][0] ;
 wire \u2.mem[47][10] ;
 wire \u2.mem[47][11] ;
 wire \u2.mem[47][12] ;
 wire \u2.mem[47][13] ;
 wire \u2.mem[47][14] ;
 wire \u2.mem[47][15] ;
 wire \u2.mem[47][1] ;
 wire \u2.mem[47][2] ;
 wire \u2.mem[47][3] ;
 wire \u2.mem[47][4] ;
 wire \u2.mem[47][5] ;
 wire \u2.mem[47][6] ;
 wire \u2.mem[47][7] ;
 wire \u2.mem[47][8] ;
 wire \u2.mem[47][9] ;
 wire \u2.mem[48][0] ;
 wire \u2.mem[48][10] ;
 wire \u2.mem[48][11] ;
 wire \u2.mem[48][12] ;
 wire \u2.mem[48][13] ;
 wire \u2.mem[48][14] ;
 wire \u2.mem[48][15] ;
 wire \u2.mem[48][1] ;
 wire \u2.mem[48][2] ;
 wire \u2.mem[48][3] ;
 wire \u2.mem[48][4] ;
 wire \u2.mem[48][5] ;
 wire \u2.mem[48][6] ;
 wire \u2.mem[48][7] ;
 wire \u2.mem[48][8] ;
 wire \u2.mem[48][9] ;
 wire \u2.mem[49][0] ;
 wire \u2.mem[49][10] ;
 wire \u2.mem[49][11] ;
 wire \u2.mem[49][12] ;
 wire \u2.mem[49][13] ;
 wire \u2.mem[49][14] ;
 wire \u2.mem[49][15] ;
 wire \u2.mem[49][1] ;
 wire \u2.mem[49][2] ;
 wire \u2.mem[49][3] ;
 wire \u2.mem[49][4] ;
 wire \u2.mem[49][5] ;
 wire \u2.mem[49][6] ;
 wire \u2.mem[49][7] ;
 wire \u2.mem[49][8] ;
 wire \u2.mem[49][9] ;
 wire \u2.mem[4][0] ;
 wire \u2.mem[4][10] ;
 wire \u2.mem[4][11] ;
 wire \u2.mem[4][12] ;
 wire \u2.mem[4][13] ;
 wire \u2.mem[4][14] ;
 wire \u2.mem[4][15] ;
 wire \u2.mem[4][1] ;
 wire \u2.mem[4][2] ;
 wire \u2.mem[4][3] ;
 wire \u2.mem[4][4] ;
 wire \u2.mem[4][5] ;
 wire \u2.mem[4][6] ;
 wire \u2.mem[4][7] ;
 wire \u2.mem[4][8] ;
 wire \u2.mem[4][9] ;
 wire \u2.mem[50][0] ;
 wire \u2.mem[50][10] ;
 wire \u2.mem[50][11] ;
 wire \u2.mem[50][12] ;
 wire \u2.mem[50][13] ;
 wire \u2.mem[50][14] ;
 wire \u2.mem[50][15] ;
 wire \u2.mem[50][1] ;
 wire \u2.mem[50][2] ;
 wire \u2.mem[50][3] ;
 wire \u2.mem[50][4] ;
 wire \u2.mem[50][5] ;
 wire \u2.mem[50][6] ;
 wire \u2.mem[50][7] ;
 wire \u2.mem[50][8] ;
 wire \u2.mem[50][9] ;
 wire \u2.mem[51][0] ;
 wire \u2.mem[51][10] ;
 wire \u2.mem[51][11] ;
 wire \u2.mem[51][12] ;
 wire \u2.mem[51][13] ;
 wire \u2.mem[51][14] ;
 wire \u2.mem[51][15] ;
 wire \u2.mem[51][1] ;
 wire \u2.mem[51][2] ;
 wire \u2.mem[51][3] ;
 wire \u2.mem[51][4] ;
 wire \u2.mem[51][5] ;
 wire \u2.mem[51][6] ;
 wire \u2.mem[51][7] ;
 wire \u2.mem[51][8] ;
 wire \u2.mem[51][9] ;
 wire \u2.mem[52][0] ;
 wire \u2.mem[52][10] ;
 wire \u2.mem[52][11] ;
 wire \u2.mem[52][12] ;
 wire \u2.mem[52][13] ;
 wire \u2.mem[52][14] ;
 wire \u2.mem[52][15] ;
 wire \u2.mem[52][1] ;
 wire \u2.mem[52][2] ;
 wire \u2.mem[52][3] ;
 wire \u2.mem[52][4] ;
 wire \u2.mem[52][5] ;
 wire \u2.mem[52][6] ;
 wire \u2.mem[52][7] ;
 wire \u2.mem[52][8] ;
 wire \u2.mem[52][9] ;
 wire \u2.mem[53][0] ;
 wire \u2.mem[53][10] ;
 wire \u2.mem[53][11] ;
 wire \u2.mem[53][12] ;
 wire \u2.mem[53][13] ;
 wire \u2.mem[53][14] ;
 wire \u2.mem[53][15] ;
 wire \u2.mem[53][1] ;
 wire \u2.mem[53][2] ;
 wire \u2.mem[53][3] ;
 wire \u2.mem[53][4] ;
 wire \u2.mem[53][5] ;
 wire \u2.mem[53][6] ;
 wire \u2.mem[53][7] ;
 wire \u2.mem[53][8] ;
 wire \u2.mem[53][9] ;
 wire \u2.mem[54][0] ;
 wire \u2.mem[54][10] ;
 wire \u2.mem[54][11] ;
 wire \u2.mem[54][12] ;
 wire \u2.mem[54][13] ;
 wire \u2.mem[54][14] ;
 wire \u2.mem[54][15] ;
 wire \u2.mem[54][1] ;
 wire \u2.mem[54][2] ;
 wire \u2.mem[54][3] ;
 wire \u2.mem[54][4] ;
 wire \u2.mem[54][5] ;
 wire \u2.mem[54][6] ;
 wire \u2.mem[54][7] ;
 wire \u2.mem[54][8] ;
 wire \u2.mem[54][9] ;
 wire \u2.mem[55][0] ;
 wire \u2.mem[55][10] ;
 wire \u2.mem[55][11] ;
 wire \u2.mem[55][12] ;
 wire \u2.mem[55][13] ;
 wire \u2.mem[55][14] ;
 wire \u2.mem[55][15] ;
 wire \u2.mem[55][1] ;
 wire \u2.mem[55][2] ;
 wire \u2.mem[55][3] ;
 wire \u2.mem[55][4] ;
 wire \u2.mem[55][5] ;
 wire \u2.mem[55][6] ;
 wire \u2.mem[55][7] ;
 wire \u2.mem[55][8] ;
 wire \u2.mem[55][9] ;
 wire \u2.mem[56][0] ;
 wire \u2.mem[56][10] ;
 wire \u2.mem[56][11] ;
 wire \u2.mem[56][12] ;
 wire \u2.mem[56][13] ;
 wire \u2.mem[56][14] ;
 wire \u2.mem[56][15] ;
 wire \u2.mem[56][1] ;
 wire \u2.mem[56][2] ;
 wire \u2.mem[56][3] ;
 wire \u2.mem[56][4] ;
 wire \u2.mem[56][5] ;
 wire \u2.mem[56][6] ;
 wire \u2.mem[56][7] ;
 wire \u2.mem[56][8] ;
 wire \u2.mem[56][9] ;
 wire \u2.mem[57][0] ;
 wire \u2.mem[57][10] ;
 wire \u2.mem[57][11] ;
 wire \u2.mem[57][12] ;
 wire \u2.mem[57][13] ;
 wire \u2.mem[57][14] ;
 wire \u2.mem[57][15] ;
 wire \u2.mem[57][1] ;
 wire \u2.mem[57][2] ;
 wire \u2.mem[57][3] ;
 wire \u2.mem[57][4] ;
 wire \u2.mem[57][5] ;
 wire \u2.mem[57][6] ;
 wire \u2.mem[57][7] ;
 wire \u2.mem[57][8] ;
 wire \u2.mem[57][9] ;
 wire \u2.mem[58][0] ;
 wire \u2.mem[58][10] ;
 wire \u2.mem[58][11] ;
 wire \u2.mem[58][12] ;
 wire \u2.mem[58][13] ;
 wire \u2.mem[58][14] ;
 wire \u2.mem[58][15] ;
 wire \u2.mem[58][1] ;
 wire \u2.mem[58][2] ;
 wire \u2.mem[58][3] ;
 wire \u2.mem[58][4] ;
 wire \u2.mem[58][5] ;
 wire \u2.mem[58][6] ;
 wire \u2.mem[58][7] ;
 wire \u2.mem[58][8] ;
 wire \u2.mem[58][9] ;
 wire \u2.mem[59][0] ;
 wire \u2.mem[59][10] ;
 wire \u2.mem[59][11] ;
 wire \u2.mem[59][12] ;
 wire \u2.mem[59][13] ;
 wire \u2.mem[59][14] ;
 wire \u2.mem[59][15] ;
 wire \u2.mem[59][1] ;
 wire \u2.mem[59][2] ;
 wire \u2.mem[59][3] ;
 wire \u2.mem[59][4] ;
 wire \u2.mem[59][5] ;
 wire \u2.mem[59][6] ;
 wire \u2.mem[59][7] ;
 wire \u2.mem[59][8] ;
 wire \u2.mem[59][9] ;
 wire \u2.mem[5][0] ;
 wire \u2.mem[5][10] ;
 wire \u2.mem[5][11] ;
 wire \u2.mem[5][12] ;
 wire \u2.mem[5][13] ;
 wire \u2.mem[5][14] ;
 wire \u2.mem[5][15] ;
 wire \u2.mem[5][1] ;
 wire \u2.mem[5][2] ;
 wire \u2.mem[5][3] ;
 wire \u2.mem[5][4] ;
 wire \u2.mem[5][5] ;
 wire \u2.mem[5][6] ;
 wire \u2.mem[5][7] ;
 wire \u2.mem[5][8] ;
 wire \u2.mem[5][9] ;
 wire \u2.mem[60][0] ;
 wire \u2.mem[60][10] ;
 wire \u2.mem[60][11] ;
 wire \u2.mem[60][12] ;
 wire \u2.mem[60][13] ;
 wire \u2.mem[60][14] ;
 wire \u2.mem[60][15] ;
 wire \u2.mem[60][1] ;
 wire \u2.mem[60][2] ;
 wire \u2.mem[60][3] ;
 wire \u2.mem[60][4] ;
 wire \u2.mem[60][5] ;
 wire \u2.mem[60][6] ;
 wire \u2.mem[60][7] ;
 wire \u2.mem[60][8] ;
 wire \u2.mem[60][9] ;
 wire \u2.mem[61][0] ;
 wire \u2.mem[61][10] ;
 wire \u2.mem[61][11] ;
 wire \u2.mem[61][12] ;
 wire \u2.mem[61][13] ;
 wire \u2.mem[61][14] ;
 wire \u2.mem[61][15] ;
 wire \u2.mem[61][1] ;
 wire \u2.mem[61][2] ;
 wire \u2.mem[61][3] ;
 wire \u2.mem[61][4] ;
 wire \u2.mem[61][5] ;
 wire \u2.mem[61][6] ;
 wire \u2.mem[61][7] ;
 wire \u2.mem[61][8] ;
 wire \u2.mem[61][9] ;
 wire \u2.mem[62][0] ;
 wire \u2.mem[62][10] ;
 wire \u2.mem[62][11] ;
 wire \u2.mem[62][12] ;
 wire \u2.mem[62][13] ;
 wire \u2.mem[62][14] ;
 wire \u2.mem[62][15] ;
 wire \u2.mem[62][1] ;
 wire \u2.mem[62][2] ;
 wire \u2.mem[62][3] ;
 wire \u2.mem[62][4] ;
 wire \u2.mem[62][5] ;
 wire \u2.mem[62][6] ;
 wire \u2.mem[62][7] ;
 wire \u2.mem[62][8] ;
 wire \u2.mem[62][9] ;
 wire \u2.mem[63][0] ;
 wire \u2.mem[63][10] ;
 wire \u2.mem[63][11] ;
 wire \u2.mem[63][12] ;
 wire \u2.mem[63][13] ;
 wire \u2.mem[63][14] ;
 wire \u2.mem[63][15] ;
 wire \u2.mem[63][1] ;
 wire \u2.mem[63][2] ;
 wire \u2.mem[63][3] ;
 wire \u2.mem[63][4] ;
 wire \u2.mem[63][5] ;
 wire \u2.mem[63][6] ;
 wire \u2.mem[63][7] ;
 wire \u2.mem[63][8] ;
 wire \u2.mem[63][9] ;
 wire \u2.mem[6][0] ;
 wire \u2.mem[6][10] ;
 wire \u2.mem[6][11] ;
 wire \u2.mem[6][12] ;
 wire \u2.mem[6][13] ;
 wire \u2.mem[6][14] ;
 wire \u2.mem[6][15] ;
 wire \u2.mem[6][1] ;
 wire \u2.mem[6][2] ;
 wire \u2.mem[6][3] ;
 wire \u2.mem[6][4] ;
 wire \u2.mem[6][5] ;
 wire \u2.mem[6][6] ;
 wire \u2.mem[6][7] ;
 wire \u2.mem[6][8] ;
 wire \u2.mem[6][9] ;
 wire \u2.mem[7][0] ;
 wire \u2.mem[7][10] ;
 wire \u2.mem[7][11] ;
 wire \u2.mem[7][12] ;
 wire \u2.mem[7][13] ;
 wire \u2.mem[7][14] ;
 wire \u2.mem[7][15] ;
 wire \u2.mem[7][1] ;
 wire \u2.mem[7][2] ;
 wire \u2.mem[7][3] ;
 wire \u2.mem[7][4] ;
 wire \u2.mem[7][5] ;
 wire \u2.mem[7][6] ;
 wire \u2.mem[7][7] ;
 wire \u2.mem[7][8] ;
 wire \u2.mem[7][9] ;
 wire \u2.mem[8][0] ;
 wire \u2.mem[8][10] ;
 wire \u2.mem[8][11] ;
 wire \u2.mem[8][12] ;
 wire \u2.mem[8][13] ;
 wire \u2.mem[8][14] ;
 wire \u2.mem[8][15] ;
 wire \u2.mem[8][1] ;
 wire \u2.mem[8][2] ;
 wire \u2.mem[8][3] ;
 wire \u2.mem[8][4] ;
 wire \u2.mem[8][5] ;
 wire \u2.mem[8][6] ;
 wire \u2.mem[8][7] ;
 wire \u2.mem[8][8] ;
 wire \u2.mem[8][9] ;
 wire \u2.mem[9][0] ;
 wire \u2.mem[9][10] ;
 wire \u2.mem[9][11] ;
 wire \u2.mem[9][12] ;
 wire \u2.mem[9][13] ;
 wire \u2.mem[9][14] ;
 wire \u2.mem[9][15] ;
 wire \u2.mem[9][1] ;
 wire \u2.mem[9][2] ;
 wire \u2.mem[9][3] ;
 wire \u2.mem[9][4] ;
 wire \u2.mem[9][5] ;
 wire \u2.mem[9][6] ;
 wire \u2.mem[9][7] ;
 wire \u2.mem[9][8] ;
 wire \u2.mem[9][9] ;
 wire \u2.select_mem_col[0] ;
 wire \u2.select_mem_col[1] ;
 wire \u2.select_mem_col[2] ;
 wire \u2.select_mem_col[3] ;
 wire \u2.select_mem_col[4] ;
 wire \u2.select_mem_col[5] ;
 wire \u2.select_mem_row[0] ;
 wire \u2.select_mem_row[1] ;
 wire \u2.select_mem_row[2] ;
 wire \u2.select_mem_row[3] ;
 wire \u2.select_mem_row[4] ;
 wire \u2.select_mem_row[5] ;
 wire \u3.data ;
 wire \u3.enable ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire clknet_leaf_0_clock;
 wire clknet_leaf_1_clock;
 wire clknet_leaf_2_clock;
 wire clknet_leaf_3_clock;
 wire clknet_leaf_4_clock;
 wire clknet_leaf_5_clock;
 wire clknet_leaf_7_clock;
 wire clknet_leaf_8_clock;
 wire clknet_leaf_9_clock;
 wire clknet_leaf_10_clock;
 wire clknet_leaf_11_clock;
 wire clknet_leaf_12_clock;
 wire clknet_leaf_13_clock;
 wire clknet_leaf_14_clock;
 wire clknet_leaf_15_clock;
 wire clknet_leaf_16_clock;
 wire clknet_leaf_17_clock;
 wire clknet_leaf_18_clock;
 wire clknet_leaf_19_clock;
 wire clknet_leaf_20_clock;
 wire clknet_leaf_21_clock;
 wire clknet_leaf_22_clock;
 wire clknet_leaf_23_clock;
 wire clknet_leaf_24_clock;
 wire clknet_leaf_25_clock;
 wire clknet_leaf_26_clock;
 wire clknet_leaf_27_clock;
 wire clknet_leaf_28_clock;
 wire clknet_leaf_29_clock;
 wire clknet_leaf_30_clock;
 wire clknet_leaf_31_clock;
 wire clknet_leaf_32_clock;
 wire clknet_leaf_33_clock;
 wire clknet_leaf_34_clock;
 wire clknet_leaf_35_clock;
 wire clknet_leaf_36_clock;
 wire clknet_leaf_37_clock;
 wire clknet_leaf_38_clock;
 wire clknet_leaf_39_clock;
 wire clknet_leaf_40_clock;
 wire clknet_leaf_41_clock;
 wire clknet_leaf_42_clock;
 wire clknet_leaf_43_clock;
 wire clknet_leaf_44_clock;
 wire clknet_leaf_45_clock;
 wire clknet_leaf_46_clock;
 wire clknet_leaf_47_clock;
 wire clknet_leaf_48_clock;
 wire clknet_leaf_49_clock;
 wire clknet_leaf_50_clock;
 wire clknet_leaf_51_clock;
 wire clknet_leaf_52_clock;
 wire clknet_leaf_53_clock;
 wire clknet_leaf_54_clock;
 wire clknet_leaf_55_clock;
 wire clknet_leaf_56_clock;
 wire clknet_leaf_57_clock;
 wire clknet_leaf_58_clock;
 wire clknet_leaf_59_clock;
 wire clknet_leaf_60_clock;
 wire clknet_leaf_61_clock;
 wire clknet_leaf_62_clock;
 wire clknet_leaf_63_clock;
 wire clknet_leaf_64_clock;
 wire clknet_leaf_65_clock;
 wire clknet_leaf_66_clock;
 wire clknet_leaf_67_clock;
 wire clknet_leaf_68_clock;
 wire clknet_leaf_69_clock;
 wire clknet_leaf_70_clock;
 wire clknet_leaf_71_clock;
 wire clknet_leaf_72_clock;
 wire clknet_leaf_73_clock;
 wire clknet_leaf_74_clock;
 wire clknet_leaf_75_clock;
 wire clknet_leaf_76_clock;
 wire clknet_leaf_77_clock;
 wire clknet_leaf_78_clock;
 wire clknet_leaf_79_clock;
 wire clknet_leaf_80_clock;
 wire clknet_leaf_81_clock;
 wire clknet_leaf_82_clock;
 wire clknet_leaf_83_clock;
 wire clknet_leaf_84_clock;
 wire clknet_leaf_85_clock;
 wire clknet_leaf_86_clock;
 wire clknet_leaf_87_clock;
 wire clknet_leaf_88_clock;
 wire clknet_leaf_89_clock;
 wire clknet_leaf_90_clock;
 wire clknet_leaf_91_clock;
 wire clknet_leaf_92_clock;
 wire clknet_leaf_93_clock;
 wire clknet_leaf_94_clock;
 wire clknet_leaf_95_clock;
 wire clknet_leaf_96_clock;
 wire clknet_leaf_97_clock;
 wire clknet_leaf_98_clock;
 wire clknet_leaf_99_clock;
 wire clknet_leaf_100_clock;
 wire clknet_leaf_101_clock;
 wire clknet_leaf_102_clock;
 wire clknet_leaf_103_clock;
 wire clknet_leaf_104_clock;
 wire clknet_leaf_105_clock;
 wire clknet_leaf_106_clock;
 wire clknet_leaf_107_clock;
 wire clknet_leaf_108_clock;
 wire clknet_leaf_109_clock;
 wire clknet_leaf_110_clock;
 wire clknet_leaf_111_clock;
 wire clknet_leaf_112_clock;
 wire clknet_leaf_113_clock;
 wire clknet_leaf_114_clock;
 wire clknet_leaf_115_clock;
 wire clknet_leaf_116_clock;
 wire clknet_leaf_117_clock;
 wire clknet_leaf_118_clock;
 wire clknet_leaf_119_clock;
 wire clknet_leaf_120_clock;
 wire clknet_leaf_121_clock;
 wire clknet_leaf_122_clock;
 wire clknet_leaf_123_clock;
 wire clknet_leaf_124_clock;
 wire clknet_leaf_125_clock;
 wire clknet_leaf_126_clock;
 wire clknet_leaf_127_clock;
 wire clknet_leaf_128_clock;
 wire clknet_leaf_129_clock;
 wire clknet_leaf_130_clock;
 wire clknet_leaf_131_clock;
 wire clknet_leaf_132_clock;
 wire clknet_leaf_133_clock;
 wire clknet_leaf_134_clock;
 wire clknet_leaf_135_clock;
 wire clknet_leaf_136_clock;
 wire clknet_leaf_137_clock;
 wire clknet_leaf_138_clock;
 wire clknet_leaf_139_clock;
 wire clknet_leaf_140_clock;
 wire clknet_leaf_141_clock;
 wire clknet_leaf_143_clock;
 wire clknet_leaf_144_clock;
 wire clknet_leaf_145_clock;
 wire clknet_leaf_146_clock;
 wire clknet_leaf_147_clock;
 wire clknet_leaf_148_clock;
 wire clknet_leaf_149_clock;
 wire clknet_leaf_150_clock;
 wire clknet_leaf_151_clock;
 wire clknet_leaf_152_clock;
 wire clknet_leaf_153_clock;
 wire clknet_leaf_154_clock;
 wire clknet_leaf_155_clock;
 wire clknet_leaf_156_clock;
 wire clknet_leaf_157_clock;
 wire clknet_leaf_158_clock;
 wire clknet_leaf_159_clock;
 wire clknet_leaf_160_clock;
 wire clknet_leaf_161_clock;
 wire clknet_leaf_162_clock;
 wire clknet_leaf_163_clock;
 wire clknet_leaf_164_clock;
 wire clknet_leaf_165_clock;
 wire clknet_leaf_166_clock;
 wire clknet_leaf_167_clock;
 wire clknet_leaf_168_clock;
 wire clknet_leaf_169_clock;
 wire clknet_leaf_170_clock;
 wire clknet_leaf_171_clock;
 wire clknet_leaf_172_clock;
 wire clknet_leaf_173_clock;
 wire clknet_leaf_174_clock;
 wire clknet_leaf_175_clock;
 wire clknet_leaf_177_clock;
 wire clknet_leaf_178_clock;
 wire clknet_leaf_179_clock;
 wire clknet_leaf_180_clock;
 wire clknet_leaf_181_clock;
 wire clknet_leaf_182_clock;
 wire clknet_leaf_183_clock;
 wire clknet_leaf_184_clock;
 wire clknet_leaf_185_clock;
 wire clknet_leaf_186_clock;
 wire clknet_leaf_187_clock;
 wire clknet_leaf_188_clock;
 wire clknet_leaf_189_clock;
 wire clknet_leaf_190_clock;
 wire clknet_leaf_191_clock;
 wire clknet_leaf_192_clock;
 wire clknet_leaf_193_clock;
 wire clknet_leaf_194_clock;
 wire clknet_leaf_195_clock;
 wire clknet_leaf_196_clock;
 wire clknet_leaf_197_clock;
 wire clknet_leaf_198_clock;
 wire clknet_leaf_199_clock;
 wire clknet_leaf_200_clock;
 wire clknet_leaf_201_clock;
 wire clknet_leaf_202_clock;
 wire clknet_leaf_203_clock;
 wire clknet_leaf_204_clock;
 wire clknet_leaf_205_clock;
 wire clknet_leaf_206_clock;
 wire clknet_leaf_207_clock;
 wire clknet_leaf_208_clock;
 wire clknet_leaf_209_clock;
 wire clknet_leaf_210_clock;
 wire clknet_leaf_211_clock;
 wire clknet_leaf_212_clock;
 wire clknet_leaf_213_clock;
 wire clknet_leaf_214_clock;
 wire clknet_leaf_215_clock;
 wire clknet_leaf_216_clock;
 wire clknet_leaf_217_clock;
 wire clknet_leaf_218_clock;
 wire clknet_leaf_219_clock;
 wire clknet_leaf_220_clock;
 wire clknet_leaf_221_clock;
 wire clknet_leaf_222_clock;
 wire clknet_leaf_223_clock;
 wire clknet_leaf_224_clock;
 wire clknet_leaf_225_clock;
 wire clknet_leaf_226_clock;
 wire clknet_leaf_227_clock;
 wire clknet_leaf_228_clock;
 wire clknet_leaf_229_clock;
 wire clknet_leaf_230_clock;
 wire clknet_leaf_231_clock;
 wire clknet_leaf_232_clock;
 wire clknet_leaf_233_clock;
 wire clknet_leaf_234_clock;
 wire clknet_leaf_235_clock;
 wire clknet_leaf_236_clock;
 wire clknet_leaf_237_clock;
 wire clknet_leaf_238_clock;
 wire clknet_leaf_239_clock;
 wire clknet_leaf_240_clock;
 wire clknet_leaf_241_clock;
 wire clknet_leaf_242_clock;
 wire clknet_leaf_243_clock;
 wire clknet_leaf_244_clock;
 wire clknet_leaf_245_clock;
 wire clknet_leaf_246_clock;
 wire clknet_leaf_248_clock;
 wire clknet_leaf_249_clock;
 wire clknet_leaf_250_clock;
 wire clknet_leaf_251_clock;
 wire clknet_leaf_252_clock;
 wire clknet_leaf_253_clock;
 wire clknet_leaf_254_clock;
 wire clknet_leaf_255_clock;
 wire clknet_leaf_256_clock;
 wire clknet_leaf_257_clock;
 wire clknet_leaf_258_clock;
 wire clknet_leaf_259_clock;
 wire clknet_leaf_260_clock;
 wire clknet_leaf_261_clock;
 wire clknet_leaf_262_clock;
 wire clknet_leaf_263_clock;
 wire clknet_leaf_264_clock;
 wire clknet_leaf_265_clock;
 wire clknet_leaf_266_clock;
 wire clknet_leaf_267_clock;
 wire clknet_leaf_268_clock;
 wire clknet_leaf_269_clock;
 wire clknet_leaf_270_clock;
 wire clknet_leaf_271_clock;
 wire clknet_leaf_272_clock;
 wire clknet_leaf_273_clock;
 wire clknet_leaf_274_clock;
 wire clknet_leaf_275_clock;
 wire clknet_leaf_276_clock;
 wire clknet_leaf_277_clock;
 wire clknet_leaf_278_clock;
 wire clknet_leaf_279_clock;
 wire clknet_leaf_280_clock;
 wire clknet_leaf_281_clock;
 wire clknet_leaf_282_clock;
 wire clknet_leaf_283_clock;
 wire clknet_leaf_284_clock;
 wire clknet_leaf_285_clock;
 wire clknet_leaf_286_clock;
 wire clknet_leaf_287_clock;
 wire clknet_leaf_288_clock;
 wire clknet_leaf_289_clock;
 wire clknet_leaf_290_clock;
 wire clknet_leaf_291_clock;
 wire clknet_leaf_292_clock;
 wire clknet_leaf_293_clock;
 wire clknet_leaf_294_clock;
 wire clknet_leaf_295_clock;
 wire clknet_leaf_296_clock;
 wire clknet_leaf_297_clock;
 wire clknet_leaf_298_clock;
 wire clknet_leaf_299_clock;
 wire clknet_leaf_300_clock;
 wire clknet_leaf_301_clock;
 wire clknet_leaf_302_clock;
 wire clknet_leaf_303_clock;
 wire clknet_leaf_304_clock;
 wire clknet_leaf_305_clock;
 wire clknet_leaf_306_clock;
 wire clknet_leaf_307_clock;
 wire clknet_leaf_309_clock;
 wire clknet_leaf_310_clock;
 wire clknet_leaf_311_clock;
 wire clknet_leaf_312_clock;
 wire clknet_leaf_313_clock;
 wire clknet_leaf_314_clock;
 wire clknet_leaf_315_clock;
 wire clknet_leaf_316_clock;
 wire clknet_leaf_317_clock;
 wire clknet_leaf_318_clock;
 wire clknet_leaf_319_clock;
 wire clknet_leaf_320_clock;
 wire clknet_leaf_321_clock;
 wire clknet_leaf_322_clock;
 wire clknet_leaf_323_clock;
 wire clknet_leaf_324_clock;
 wire clknet_leaf_325_clock;
 wire clknet_leaf_326_clock;
 wire clknet_leaf_327_clock;
 wire clknet_leaf_328_clock;
 wire clknet_leaf_329_clock;
 wire clknet_leaf_330_clock;
 wire clknet_leaf_331_clock;
 wire clknet_leaf_332_clock;
 wire clknet_leaf_333_clock;
 wire clknet_leaf_334_clock;
 wire clknet_leaf_335_clock;
 wire clknet_leaf_336_clock;
 wire clknet_leaf_337_clock;
 wire clknet_leaf_338_clock;
 wire clknet_leaf_340_clock;
 wire clknet_leaf_341_clock;
 wire clknet_leaf_342_clock;
 wire clknet_leaf_343_clock;
 wire clknet_leaf_344_clock;
 wire clknet_leaf_345_clock;
 wire clknet_leaf_346_clock;
 wire clknet_leaf_347_clock;
 wire clknet_leaf_348_clock;
 wire clknet_leaf_349_clock;
 wire clknet_leaf_350_clock;
 wire clknet_leaf_352_clock;
 wire clknet_leaf_353_clock;
 wire clknet_leaf_354_clock;
 wire clknet_leaf_355_clock;
 wire clknet_leaf_356_clock;
 wire clknet_leaf_357_clock;
 wire clknet_leaf_358_clock;
 wire clknet_leaf_359_clock;
 wire clknet_leaf_360_clock;
 wire clknet_leaf_361_clock;
 wire clknet_leaf_362_clock;
 wire clknet_leaf_363_clock;
 wire clknet_leaf_364_clock;
 wire clknet_0_clock;
 wire clknet_3_0_0_clock;
 wire clknet_3_1_0_clock;
 wire clknet_3_2_0_clock;
 wire clknet_3_3_0_clock;
 wire clknet_3_4_0_clock;
 wire clknet_3_5_0_clock;
 wire clknet_3_6_0_clock;
 wire clknet_3_7_0_clock;
 wire clknet_4_0_0_clock;
 wire clknet_4_1_0_clock;
 wire clknet_4_2_0_clock;
 wire clknet_4_3_0_clock;
 wire clknet_4_4_0_clock;
 wire clknet_4_5_0_clock;
 wire clknet_4_6_0_clock;
 wire clknet_4_7_0_clock;
 wire clknet_4_8_0_clock;
 wire clknet_4_9_0_clock;
 wire clknet_4_10_0_clock;
 wire clknet_4_11_0_clock;
 wire clknet_4_12_0_clock;
 wire clknet_4_13_0_clock;
 wire clknet_4_14_0_clock;
 wire clknet_4_15_0_clock;
 wire clknet_5_0_0_clock;
 wire clknet_5_1_0_clock;
 wire clknet_5_2_0_clock;
 wire clknet_5_3_0_clock;
 wire clknet_5_4_0_clock;
 wire clknet_5_5_0_clock;
 wire clknet_5_6_0_clock;
 wire clknet_5_7_0_clock;
 wire clknet_5_8_0_clock;
 wire clknet_5_9_0_clock;
 wire clknet_5_10_0_clock;
 wire clknet_5_11_0_clock;
 wire clknet_5_12_0_clock;
 wire clknet_5_13_0_clock;
 wire clknet_5_14_0_clock;
 wire clknet_5_15_0_clock;
 wire clknet_5_16_0_clock;
 wire clknet_5_17_0_clock;
 wire clknet_5_18_0_clock;
 wire clknet_5_19_0_clock;
 wire clknet_5_20_0_clock;
 wire clknet_5_21_0_clock;
 wire clknet_5_22_0_clock;
 wire clknet_5_23_0_clock;
 wire clknet_5_24_0_clock;
 wire clknet_5_25_0_clock;
 wire clknet_5_26_0_clock;
 wire clknet_5_27_0_clock;
 wire clknet_5_28_0_clock;
 wire clknet_5_29_0_clock;
 wire clknet_5_30_0_clock;
 wire clknet_5_31_0_clock;
 wire clknet_0_clock_a;
 wire clknet_2_0__leaf_clock_a;
 wire clknet_2_1__leaf_clock_a;
 wire clknet_2_2__leaf_clock_a;
 wire clknet_2_3__leaf_clock_a;
 wire net45;

 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05993_ (.I(\row_col_select_trans.data_sync ),
    .Z(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05994_ (.I0(\u2.select_mem_row[1] ),
    .I1(\u2.select_mem_col[1] ),
    .S(_01502_),
    .Z(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05995_ (.I(_01503_),
    .Z(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05996_ (.I(\u2.select_mem_col[0] ),
    .ZN(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05997_ (.A1(\u2.select_mem_row[0] ),
    .A2(\row_col_select_trans.data_sync ),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05998_ (.A1(_01505_),
    .A2(\row_col_select_trans.data_sync ),
    .B(_01506_),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05999_ (.I(_01507_),
    .Z(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06000_ (.A1(\u2.driver_mem[3] ),
    .A2(_01508_),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06001_ (.I(_01502_),
    .Z(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06002_ (.A1(_01505_),
    .A2(_01502_),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06003_ (.A1(\u2.select_mem_row[0] ),
    .A2(_01510_),
    .B(_01511_),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06004_ (.I(_01512_),
    .Z(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06005_ (.A1(\u2.driver_mem[2] ),
    .A2(_01513_),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06006_ (.A1(_01504_),
    .A2(_01509_),
    .A3(_01514_),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06007_ (.I0(\u2.select_mem_row[2] ),
    .I1(\u2.select_mem_col[2] ),
    .S(_01510_),
    .Z(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06008_ (.I(_01512_),
    .Z(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06009_ (.I(_01507_),
    .Z(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06010_ (.A1(\u2.driver_mem[1] ),
    .A2(_01518_),
    .Z(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06011_ (.I(_01503_),
    .Z(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06012_ (.A1(\u2.driver_mem[0] ),
    .A2(_01517_),
    .B(_01519_),
    .C(_01520_),
    .ZN(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06013_ (.A1(_01516_),
    .A2(_01521_),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06014_ (.A1(\u2.driver_mem[7] ),
    .A2(_01508_),
    .Z(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06015_ (.A1(\u2.driver_mem[6] ),
    .A2(_01513_),
    .B(_01523_),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06016_ (.A1(\u2.driver_mem[5] ),
    .A2(_01518_),
    .Z(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06017_ (.A1(\u2.driver_mem[4] ),
    .A2(_01517_),
    .B(_01525_),
    .C(_01520_),
    .ZN(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06018_ (.A1(_01504_),
    .A2(_01524_),
    .B(_01526_),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06019_ (.A1(_01515_),
    .A2(_01522_),
    .B1(_01527_),
    .B2(_01516_),
    .ZN(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06020_ (.A1(\u2.driver_mem[11] ),
    .A2(_01508_),
    .ZN(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06021_ (.A1(\u2.driver_mem[10] ),
    .A2(_01513_),
    .ZN(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06022_ (.A1(_01504_),
    .A2(_01529_),
    .A3(_01530_),
    .ZN(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06023_ (.A1(\u2.driver_mem[9] ),
    .A2(_01518_),
    .Z(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06024_ (.A1(\u2.driver_mem[8] ),
    .A2(_01517_),
    .B(_01532_),
    .C(_01520_),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06025_ (.A1(_01516_),
    .A2(_01533_),
    .ZN(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06026_ (.A1(\u2.driver_mem[15] ),
    .A2(_01508_),
    .Z(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06027_ (.A1(\u2.driver_mem[14] ),
    .A2(_01513_),
    .B(_01535_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06028_ (.A1(\u2.driver_mem[13] ),
    .A2(_01518_),
    .Z(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06029_ (.A1(\u2.driver_mem[12] ),
    .A2(_01517_),
    .B(_01537_),
    .C(_01520_),
    .ZN(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06030_ (.A1(_01504_),
    .A2(_01536_),
    .B(_01538_),
    .ZN(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06031_ (.A1(_01531_),
    .A2(_01534_),
    .B1(_01539_),
    .B2(_01516_),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06032_ (.I0(\u2.select_mem_row[3] ),
    .I1(\u2.select_mem_col[3] ),
    .S(_01510_),
    .Z(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06033_ (.I0(_01528_),
    .I1(_01540_),
    .S(_01541_),
    .Z(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06034_ (.A1(\inverter_select_trans.data_sync ),
    .A2(_01542_),
    .ZN(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06035_ (.I(_01543_),
    .Z(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06036_ (.A1(\u3.data ),
    .A2(\u3.enable ),
    .ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06037_ (.I(\u2.mem[0][0] ),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06038_ (.I(_01544_),
    .Z(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06039_ (.A1(\col_select_trans[0].data_sync ),
    .A2(\col_select_trans[1].data_sync ),
    .ZN(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06040_ (.I(_01546_),
    .Z(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06041_ (.A1(\col_select_trans[2].data_sync ),
    .A2(\col_select_trans[3].data_sync ),
    .ZN(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06042_ (.I(_01548_),
    .Z(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06043_ (.I(\col_select_trans[5].data_sync ),
    .Z(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06044_ (.I(\col_select_trans[4].data_sync ),
    .Z(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06045_ (.A1(_01550_),
    .A2(_01551_),
    .ZN(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06046_ (.A1(_01547_),
    .A2(_01549_),
    .B(_01552_),
    .ZN(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06047_ (.I(_01553_),
    .Z(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06048_ (.I(_01554_),
    .Z(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06049_ (.A1(_01550_),
    .A2(_01551_),
    .Z(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06050_ (.I(_01556_),
    .Z(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06051_ (.I(\col_select_trans[2].data_sync ),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06052_ (.I(\col_select_trans[3].data_sync ),
    .Z(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06053_ (.A1(_01558_),
    .A2(_01559_),
    .ZN(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06054_ (.I(_01560_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06055_ (.I(\col_select_trans[0].data_sync ),
    .ZN(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06056_ (.A1(_01562_),
    .A2(\col_select_trans[1].data_sync ),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06057_ (.I(_01563_),
    .Z(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06058_ (.A1(_01557_),
    .A2(_01561_),
    .A3(_01564_),
    .ZN(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06059_ (.I(_01556_),
    .Z(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06060_ (.I(_01566_),
    .Z(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06061_ (.I(\col_select_trans[3].data_sync ),
    .ZN(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06062_ (.A1(_01558_),
    .A2(_01568_),
    .ZN(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06063_ (.I(_01569_),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06064_ (.A1(_01547_),
    .A2(_01570_),
    .Z(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06065_ (.A1(_01567_),
    .A2(_01571_),
    .ZN(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06066_ (.I(\col_select_trans[0].data_sync ),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06067_ (.I(\col_select_trans[1].data_sync ),
    .Z(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06068_ (.I(_01574_),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06069_ (.A1(_01573_),
    .A2(_01575_),
    .A3(_01549_),
    .ZN(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06070_ (.A1(_01552_),
    .A2(_01576_),
    .ZN(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06071_ (.A1(\u2.mem[158][0] ),
    .A2(_01565_),
    .B1(_01572_),
    .B2(\u2.mem[151][0] ),
    .C1(_01577_),
    .C2(\u2.mem[193][0] ),
    .ZN(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06072_ (.I(_01551_),
    .ZN(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06073_ (.A1(_01550_),
    .A2(_01579_),
    .ZN(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06074_ (.I(_01580_),
    .Z(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06075_ (.I(_01581_),
    .Z(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06076_ (.A1(_01582_),
    .A2(_01576_),
    .ZN(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06077_ (.I(\col_select_trans[2].data_sync ),
    .ZN(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06078_ (.A1(_01573_),
    .A2(_01574_),
    .ZN(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06079_ (.A1(_01584_),
    .A2(_01559_),
    .A3(_01585_),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06080_ (.A1(_01550_),
    .A2(_01579_),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06081_ (.I(_01587_),
    .Z(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06082_ (.A1(_01586_),
    .A2(_01588_),
    .ZN(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06083_ (.A1(\u2.mem[177][0] ),
    .A2(_01583_),
    .B1(_01589_),
    .B2(\u2.mem[168][0] ),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06084_ (.I(_01570_),
    .Z(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06085_ (.A1(_01564_),
    .A2(_01591_),
    .A3(_01588_),
    .ZN(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06086_ (.A1(_01573_),
    .A2(_01575_),
    .ZN(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06087_ (.A1(_01556_),
    .A2(_01569_),
    .A3(_01593_),
    .ZN(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06088_ (.I(_01594_),
    .Z(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06089_ (.I(_01587_),
    .Z(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06090_ (.A1(_01576_),
    .A2(_01596_),
    .ZN(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06091_ (.A1(\u2.mem[166][0] ),
    .A2(_01592_),
    .B1(_01595_),
    .B2(\u2.mem[149][0] ),
    .C1(_01597_),
    .C2(\u2.mem[161][0] ),
    .ZN(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06092_ (.A1(_01546_),
    .A2(_01560_),
    .Z(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06093_ (.I(_01587_),
    .Z(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06094_ (.A1(_01599_),
    .A2(_01600_),
    .ZN(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06095_ (.I(_01601_),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06096_ (.A1(_01566_),
    .A2(_01599_),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06097_ (.I(_01603_),
    .Z(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06098_ (.A1(\u2.mem[175][0] ),
    .A2(_01602_),
    .B1(_01604_),
    .B2(\u2.mem[159][0] ),
    .ZN(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06099_ (.A1(_01578_),
    .A2(_01590_),
    .A3(_01598_),
    .A4(_01605_),
    .Z(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06100_ (.I(_01600_),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06101_ (.A1(_01584_),
    .A2(_01559_),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06102_ (.A1(_01547_),
    .A2(_01608_),
    .Z(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06103_ (.A1(_01607_),
    .A2(_01609_),
    .ZN(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06104_ (.I(_01610_),
    .Z(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06105_ (.I(_01561_),
    .Z(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06106_ (.I(_01593_),
    .Z(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06107_ (.A1(_01567_),
    .A2(_01612_),
    .A3(_01613_),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06108_ (.A1(_01562_),
    .A2(_01574_),
    .A3(_01548_),
    .ZN(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06109_ (.I(_01580_),
    .Z(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06110_ (.I(_01616_),
    .Z(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06111_ (.A1(_01615_),
    .A2(_01617_),
    .ZN(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06112_ (.A1(_01558_),
    .A2(_01568_),
    .A3(_01585_),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06113_ (.A1(_01619_),
    .A2(_01607_),
    .ZN(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06114_ (.A1(\u2.mem[178][0] ),
    .A2(_01618_),
    .B1(_01620_),
    .B2(\u2.mem[164][0] ),
    .ZN(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06115_ (.A1(_01571_),
    .A2(_01607_),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06116_ (.A1(_01571_),
    .A2(_01617_),
    .ZN(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06117_ (.A1(\u2.mem[167][0] ),
    .A2(_01622_),
    .B1(_01623_),
    .B2(\u2.mem[183][0] ),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06118_ (.A1(_01586_),
    .A2(_01617_),
    .ZN(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06119_ (.A1(\u2.mem[184][0] ),
    .A2(_01625_),
    .B(_01553_),
    .ZN(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06120_ (.A1(_01621_),
    .A2(_01624_),
    .A3(_01626_),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06121_ (.A1(\u2.mem[171][0] ),
    .A2(_01611_),
    .B1(_01614_),
    .B2(\u2.mem[157][0] ),
    .C(_01627_),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06122_ (.A1(_01558_),
    .A2(_01559_),
    .A3(_01585_),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06123_ (.A1(_01581_),
    .A2(_01629_),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06124_ (.I(_01630_),
    .Z(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06125_ (.A1(_01616_),
    .A2(_01609_),
    .ZN(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06126_ (.I(_01632_),
    .Z(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06127_ (.A1(_01549_),
    .A2(_01585_),
    .ZN(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06128_ (.A1(_01552_),
    .A2(_01634_),
    .ZN(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06129_ (.I(_01635_),
    .Z(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06130_ (.A1(\u2.mem[188][0] ),
    .A2(_01631_),
    .B1(_01633_),
    .B2(\u2.mem[187][0] ),
    .C1(_01636_),
    .C2(\u2.mem[192][0] ),
    .ZN(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06131_ (.I(_01557_),
    .Z(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06132_ (.A1(_01638_),
    .A2(_01576_),
    .ZN(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06133_ (.I(_01639_),
    .Z(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06134_ (.A1(_01573_),
    .A2(_01574_),
    .A3(_01548_),
    .ZN(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06135_ (.A1(_01641_),
    .A2(_01596_),
    .ZN(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06136_ (.I(_01642_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06137_ (.I(_01593_),
    .Z(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06138_ (.A1(_01570_),
    .A2(_01644_),
    .A3(_01600_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06139_ (.I(_01645_),
    .Z(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06140_ (.A1(\u2.mem[145][0] ),
    .A2(_01640_),
    .B1(_01643_),
    .B2(\u2.mem[163][0] ),
    .C1(\u2.mem[165][0] ),
    .C2(_01646_),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06141_ (.A1(_01606_),
    .A2(_01628_),
    .A3(_01637_),
    .A4(_01647_),
    .ZN(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06142_ (.A1(_01612_),
    .A2(_01616_),
    .A3(_01644_),
    .ZN(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06143_ (.I(_01649_),
    .Z(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06144_ (.A1(_01582_),
    .A2(_01634_),
    .ZN(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06145_ (.I(_01651_),
    .Z(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06146_ (.A1(_01607_),
    .A2(_01629_),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06147_ (.I(_01653_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06148_ (.A1(\u2.mem[189][0] ),
    .A2(_01650_),
    .B1(_01652_),
    .B2(\u2.mem[176][0] ),
    .C1(\u2.mem[172][0] ),
    .C2(_01654_),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06149_ (.A1(_01561_),
    .A2(_01564_),
    .A3(_01588_),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06150_ (.I(_01656_),
    .Z(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06151_ (.A1(_01567_),
    .A2(_01609_),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06152_ (.I(_01658_),
    .Z(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06153_ (.A1(_01570_),
    .A2(_01616_),
    .A3(_01644_),
    .ZN(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06154_ (.I(_01660_),
    .Z(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06155_ (.A1(\u2.mem[174][0] ),
    .A2(_01657_),
    .B1(_01659_),
    .B2(\u2.mem[155][0] ),
    .C1(_01661_),
    .C2(\u2.mem[181][0] ),
    .ZN(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06156_ (.A1(_01617_),
    .A2(_01619_),
    .ZN(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06157_ (.I(_01663_),
    .Z(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06158_ (.I(_01564_),
    .Z(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06159_ (.A1(_01638_),
    .A2(_01665_),
    .A3(_01591_),
    .ZN(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06160_ (.I(_01666_),
    .Z(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06161_ (.A1(\u2.mem[180][0] ),
    .A2(_01664_),
    .B1(_01667_),
    .B2(\u2.mem[150][0] ),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06162_ (.A1(_01655_),
    .A2(_01662_),
    .A3(_01668_),
    .ZN(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06163_ (.A1(_01638_),
    .A2(_01634_),
    .ZN(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06164_ (.I(_01670_),
    .Z(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06165_ (.A1(_01665_),
    .A2(_01591_),
    .A3(_01582_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06166_ (.I(_01672_),
    .Z(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06167_ (.A1(\u2.mem[144][0] ),
    .A2(_01671_),
    .B1(_01673_),
    .B2(\u2.mem[182][0] ),
    .ZN(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06168_ (.A1(_01638_),
    .A2(_01641_),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06169_ (.I(_01675_),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06170_ (.I(_01608_),
    .Z(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06171_ (.I(_01677_),
    .Z(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06172_ (.A1(_01678_),
    .A2(_01644_),
    .A3(_01588_),
    .ZN(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06173_ (.I(_01679_),
    .Z(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06174_ (.A1(_01581_),
    .A2(_01599_),
    .ZN(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06175_ (.I(_01681_),
    .Z(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06176_ (.A1(_01581_),
    .A2(_01641_),
    .ZN(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06177_ (.I(_01683_),
    .Z(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06178_ (.A1(\u2.mem[191][0] ),
    .A2(_01682_),
    .B1(_01684_),
    .B2(\u2.mem[179][0] ),
    .ZN(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06179_ (.A1(_01563_),
    .A2(_01677_),
    .A3(_01587_),
    .ZN(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06180_ (.I(_01686_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06181_ (.A1(_01566_),
    .A2(_01629_),
    .ZN(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06182_ (.I(_01688_),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06183_ (.A1(\u2.mem[170][0] ),
    .A2(_01687_),
    .B1(_01689_),
    .B2(\u2.mem[156][0] ),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06184_ (.A1(_01566_),
    .A2(_01615_),
    .ZN(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06185_ (.I(_01691_),
    .Z(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06186_ (.A1(_01563_),
    .A2(_01677_),
    .A3(_01580_),
    .ZN(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06187_ (.I(_01693_),
    .Z(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06188_ (.A1(\u2.mem[146][0] ),
    .A2(_01692_),
    .B1(_01694_),
    .B2(\u2.mem[186][0] ),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06189_ (.A1(_01685_),
    .A2(_01690_),
    .A3(_01695_),
    .ZN(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06190_ (.A1(\u2.mem[147][0] ),
    .A2(_01676_),
    .B1(_01680_),
    .B2(\u2.mem[169][0] ),
    .C(_01696_),
    .ZN(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06191_ (.A1(_01567_),
    .A2(_01665_),
    .A3(_01678_),
    .ZN(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06192_ (.I(_01698_),
    .Z(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06193_ (.A1(_01615_),
    .A2(_01596_),
    .ZN(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06194_ (.I(_01700_),
    .Z(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06195_ (.A1(_01561_),
    .A2(_01563_),
    .A3(_01580_),
    .ZN(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06196_ (.I(_01702_),
    .Z(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06197_ (.A1(_01552_),
    .A2(_01615_),
    .ZN(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06198_ (.I(_01704_),
    .Z(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06199_ (.A1(\u2.mem[190][0] ),
    .A2(_01703_),
    .B1(_01705_),
    .B2(\u2.mem[194][0] ),
    .ZN(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06200_ (.A1(_01556_),
    .A2(_01677_),
    .A3(_01593_),
    .ZN(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06201_ (.I(_01707_),
    .Z(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06202_ (.A1(_01600_),
    .A2(_01634_),
    .ZN(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06203_ (.I(_01709_),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06204_ (.A1(\u2.mem[153][0] ),
    .A2(_01708_),
    .B1(_01710_),
    .B2(\u2.mem[160][0] ),
    .ZN(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06205_ (.A1(_01557_),
    .A2(_01586_),
    .ZN(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06206_ (.I(_01712_),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06207_ (.A1(_01557_),
    .A2(_01619_),
    .ZN(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06208_ (.I(_01714_),
    .Z(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06209_ (.A1(\u2.mem[152][0] ),
    .A2(_01713_),
    .B1(_01715_),
    .B2(\u2.mem[148][0] ),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06210_ (.A1(_01706_),
    .A2(_01711_),
    .A3(_01716_),
    .ZN(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06211_ (.A1(\u2.mem[154][0] ),
    .A2(_01699_),
    .B1(_01701_),
    .B2(\u2.mem[162][0] ),
    .C(_01717_),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06212_ (.A1(_01612_),
    .A2(_01613_),
    .A3(_01596_),
    .ZN(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06213_ (.I(_01719_),
    .Z(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06214_ (.A1(_01678_),
    .A2(_01582_),
    .A3(_01613_),
    .ZN(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06215_ (.I(_01721_),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06216_ (.A1(\u2.mem[173][0] ),
    .A2(_01720_),
    .B1(_01722_),
    .B2(\u2.mem[185][0] ),
    .ZN(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06217_ (.A1(_01674_),
    .A2(_01697_),
    .A3(_01718_),
    .A4(_01723_),
    .ZN(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06218_ (.A1(_01648_),
    .A2(_01669_),
    .A3(_01724_),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06219_ (.A1(_01545_),
    .A2(_01555_),
    .B(_01725_),
    .ZN(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06220_ (.I(\u2.mem[0][1] ),
    .ZN(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06221_ (.I(_01726_),
    .Z(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06222_ (.I(_01565_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06223_ (.I(_01572_),
    .Z(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06224_ (.A1(\u2.mem[163][1] ),
    .A2(_01643_),
    .B1(_01646_),
    .B2(\u2.mem[165][1] ),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06225_ (.I(_01577_),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06226_ (.I(_01589_),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06227_ (.A1(\u2.mem[193][1] ),
    .A2(_01731_),
    .B1(_01732_),
    .B2(\u2.mem[168][1] ),
    .ZN(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06228_ (.I(_01583_),
    .Z(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06229_ (.A1(\u2.mem[145][1] ),
    .A2(_01640_),
    .B1(_01734_),
    .B2(\u2.mem[177][1] ),
    .ZN(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06230_ (.A1(_01730_),
    .A2(_01733_),
    .A3(_01735_),
    .ZN(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06231_ (.A1(\u2.mem[158][1] ),
    .A2(_01728_),
    .B1(_01729_),
    .B2(\u2.mem[151][1] ),
    .C(_01736_),
    .ZN(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06232_ (.A1(\u2.mem[144][1] ),
    .A2(_01671_),
    .B1(_01673_),
    .B2(\u2.mem[182][1] ),
    .ZN(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06233_ (.A1(\u2.mem[173][1] ),
    .A2(_01720_),
    .B1(_01722_),
    .B2(\u2.mem[185][1] ),
    .ZN(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06234_ (.A1(\u2.mem[170][1] ),
    .A2(_01687_),
    .B1(_01689_),
    .B2(\u2.mem[156][1] ),
    .ZN(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06235_ (.A1(\u2.mem[191][1] ),
    .A2(_01682_),
    .B1(_01684_),
    .B2(\u2.mem[179][1] ),
    .ZN(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06236_ (.A1(\u2.mem[146][1] ),
    .A2(_01692_),
    .B1(_01694_),
    .B2(\u2.mem[186][1] ),
    .ZN(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06237_ (.A1(_01740_),
    .A2(_01741_),
    .A3(_01742_),
    .ZN(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06238_ (.A1(\u2.mem[147][1] ),
    .A2(_01676_),
    .B1(_01680_),
    .B2(\u2.mem[169][1] ),
    .C(_01743_),
    .ZN(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06239_ (.A1(_01738_),
    .A2(_01739_),
    .A3(_01744_),
    .ZN(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06240_ (.A1(\u2.mem[178][1] ),
    .A2(_01618_),
    .B1(_01620_),
    .B2(\u2.mem[164][1] ),
    .ZN(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06241_ (.A1(\u2.mem[167][1] ),
    .A2(_01622_),
    .B1(_01623_),
    .B2(\u2.mem[183][1] ),
    .ZN(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06242_ (.A1(\u2.mem[171][1] ),
    .A2(_01610_),
    .B1(_01614_),
    .B2(\u2.mem[157][1] ),
    .ZN(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06243_ (.I(_01553_),
    .Z(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06244_ (.A1(\u2.mem[184][1] ),
    .A2(_01625_),
    .B(_01749_),
    .ZN(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06245_ (.A1(_01746_),
    .A2(_01747_),
    .A3(_01748_),
    .A4(_01750_),
    .ZN(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06246_ (.A1(\u2.mem[159][1] ),
    .A2(_01604_),
    .B1(_01595_),
    .B2(\u2.mem[149][1] ),
    .ZN(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06247_ (.I(_01592_),
    .Z(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06248_ (.I(_01597_),
    .Z(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06249_ (.A1(\u2.mem[166][1] ),
    .A2(_01753_),
    .B1(_01754_),
    .B2(\u2.mem[161][1] ),
    .ZN(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06250_ (.A1(\u2.mem[187][1] ),
    .A2(_01633_),
    .B1(_01636_),
    .B2(\u2.mem[192][1] ),
    .ZN(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06251_ (.A1(\u2.mem[175][1] ),
    .A2(_01602_),
    .B1(_01631_),
    .B2(\u2.mem[188][1] ),
    .ZN(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06252_ (.A1(_01752_),
    .A2(_01755_),
    .A3(_01756_),
    .A4(_01757_),
    .ZN(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06253_ (.A1(\u2.mem[174][1] ),
    .A2(_01656_),
    .B1(_01658_),
    .B2(\u2.mem[155][1] ),
    .C1(_01660_),
    .C2(\u2.mem[181][1] ),
    .ZN(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06254_ (.A1(\u2.mem[180][1] ),
    .A2(_01664_),
    .B1(_01666_),
    .B2(\u2.mem[150][1] ),
    .ZN(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06255_ (.A1(\u2.mem[152][1] ),
    .A2(_01713_),
    .B1(_01708_),
    .B2(\u2.mem[153][1] ),
    .ZN(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06256_ (.A1(\u2.mem[148][1] ),
    .A2(_01715_),
    .B1(_01698_),
    .B2(\u2.mem[154][1] ),
    .C1(\u2.mem[162][1] ),
    .C2(_01700_),
    .ZN(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06257_ (.A1(\u2.mem[190][1] ),
    .A2(_01703_),
    .B1(_01710_),
    .B2(\u2.mem[160][1] ),
    .C1(_01705_),
    .C2(\u2.mem[194][1] ),
    .ZN(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06258_ (.A1(\u2.mem[189][1] ),
    .A2(_01649_),
    .B1(_01651_),
    .B2(\u2.mem[176][1] ),
    .C1(\u2.mem[172][1] ),
    .C2(_01653_),
    .ZN(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06259_ (.A1(_01761_),
    .A2(_01762_),
    .A3(_01763_),
    .A4(_01764_),
    .Z(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06260_ (.A1(_01759_),
    .A2(_01760_),
    .A3(_01765_),
    .ZN(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06261_ (.A1(_01745_),
    .A2(_01751_),
    .A3(_01758_),
    .A4(_01766_),
    .ZN(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06262_ (.A1(_01727_),
    .A2(_01554_),
    .B1(_01737_),
    .B2(_01767_),
    .ZN(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06263_ (.I(\u2.mem[0][2] ),
    .ZN(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06264_ (.I(_01768_),
    .Z(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06265_ (.I(_01614_),
    .Z(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06266_ (.A1(\u2.mem[171][2] ),
    .A2(_01611_),
    .B1(_01770_),
    .B2(\u2.mem[157][2] ),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06267_ (.I(_01618_),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06268_ (.I(_01620_),
    .Z(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06269_ (.A1(\u2.mem[178][2] ),
    .A2(_01772_),
    .B1(_01773_),
    .B2(\u2.mem[164][2] ),
    .ZN(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06270_ (.I(_01622_),
    .Z(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06271_ (.I(_01623_),
    .Z(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06272_ (.A1(\u2.mem[167][2] ),
    .A2(_01775_),
    .B1(_01776_),
    .B2(\u2.mem[183][2] ),
    .ZN(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06273_ (.I(_01625_),
    .Z(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06274_ (.A1(\u2.mem[184][2] ),
    .A2(_01778_),
    .B(_01554_),
    .ZN(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06275_ (.A1(_01771_),
    .A2(_01774_),
    .A3(_01777_),
    .A4(_01779_),
    .ZN(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06276_ (.A1(\u2.mem[189][2] ),
    .A2(_01649_),
    .B1(_01663_),
    .B2(\u2.mem[180][2] ),
    .C1(_01651_),
    .C2(\u2.mem[176][2] ),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06277_ (.A1(\u2.mem[174][2] ),
    .A2(_01657_),
    .B1(_01658_),
    .B2(\u2.mem[155][2] ),
    .C1(_01661_),
    .C2(\u2.mem[181][2] ),
    .ZN(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06278_ (.A1(\u2.mem[172][2] ),
    .A2(_01654_),
    .B1(_01667_),
    .B2(\u2.mem[150][2] ),
    .ZN(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06279_ (.A1(_01781_),
    .A2(_01782_),
    .A3(_01783_),
    .ZN(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06280_ (.A1(\u2.mem[187][2] ),
    .A2(_01633_),
    .B1(_01636_),
    .B2(\u2.mem[192][2] ),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06281_ (.A1(\u2.mem[175][2] ),
    .A2(_01602_),
    .B1(_01631_),
    .B2(\u2.mem[188][2] ),
    .ZN(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06282_ (.A1(\u2.mem[159][2] ),
    .A2(_01604_),
    .B1(_01595_),
    .B2(\u2.mem[149][2] ),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06283_ (.A1(_01785_),
    .A2(_01786_),
    .A3(_01787_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06284_ (.A1(\u2.mem[166][2] ),
    .A2(_01753_),
    .B1(_01754_),
    .B2(\u2.mem[161][2] ),
    .C(_01788_),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06285_ (.A1(\u2.mem[145][2] ),
    .A2(_01639_),
    .B1(_01643_),
    .B2(\u2.mem[163][2] ),
    .C1(\u2.mem[165][2] ),
    .C2(_01645_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06286_ (.A1(\u2.mem[158][2] ),
    .A2(_01565_),
    .B1(_01572_),
    .B2(\u2.mem[151][2] ),
    .C1(_01589_),
    .C2(\u2.mem[168][2] ),
    .ZN(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06287_ (.A1(\u2.mem[193][2] ),
    .A2(_01731_),
    .B1(_01734_),
    .B2(\u2.mem[177][2] ),
    .ZN(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06288_ (.A1(_01789_),
    .A2(_01790_),
    .A3(_01791_),
    .A4(_01792_),
    .ZN(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06289_ (.A1(\u2.mem[190][2] ),
    .A2(_01703_),
    .B1(_01705_),
    .B2(\u2.mem[194][2] ),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06290_ (.A1(\u2.mem[153][2] ),
    .A2(_01708_),
    .B1(_01710_),
    .B2(\u2.mem[160][2] ),
    .ZN(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06291_ (.A1(\u2.mem[152][2] ),
    .A2(_01713_),
    .B1(_01715_),
    .B2(\u2.mem[148][2] ),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06292_ (.A1(_01794_),
    .A2(_01795_),
    .A3(_01796_),
    .ZN(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06293_ (.A1(\u2.mem[154][2] ),
    .A2(_01699_),
    .B1(_01701_),
    .B2(\u2.mem[162][2] ),
    .C(_01797_),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06294_ (.A1(\u2.mem[144][2] ),
    .A2(_01671_),
    .B1(_01673_),
    .B2(\u2.mem[182][2] ),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06295_ (.A1(\u2.mem[173][2] ),
    .A2(_01720_),
    .B1(_01722_),
    .B2(\u2.mem[185][2] ),
    .ZN(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06296_ (.A1(\u2.mem[170][2] ),
    .A2(_01687_),
    .B1(_01689_),
    .B2(\u2.mem[156][2] ),
    .ZN(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06297_ (.A1(\u2.mem[191][2] ),
    .A2(_01682_),
    .B1(_01684_),
    .B2(\u2.mem[179][2] ),
    .ZN(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06298_ (.A1(\u2.mem[146][2] ),
    .A2(_01692_),
    .B1(_01694_),
    .B2(\u2.mem[186][2] ),
    .ZN(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06299_ (.A1(_01801_),
    .A2(_01802_),
    .A3(_01803_),
    .ZN(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06300_ (.A1(\u2.mem[147][2] ),
    .A2(_01676_),
    .B1(_01680_),
    .B2(\u2.mem[169][2] ),
    .C(_01804_),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06301_ (.A1(_01798_),
    .A2(_01799_),
    .A3(_01800_),
    .A4(_01805_),
    .ZN(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06302_ (.A1(_01780_),
    .A2(_01784_),
    .A3(_01793_),
    .A4(_01806_),
    .ZN(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06303_ (.A1(_01769_),
    .A2(_01555_),
    .B(_01807_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06304_ (.I(\u2.mem[0][3] ),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06305_ (.I(_01808_),
    .Z(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06306_ (.A1(\u2.mem[178][3] ),
    .A2(_01772_),
    .B1(_01773_),
    .B2(\u2.mem[164][3] ),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06307_ (.A1(\u2.mem[167][3] ),
    .A2(_01775_),
    .B1(_01776_),
    .B2(\u2.mem[183][3] ),
    .ZN(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06308_ (.A1(\u2.mem[171][3] ),
    .A2(_01611_),
    .B1(_01770_),
    .B2(\u2.mem[157][3] ),
    .ZN(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06309_ (.A1(\u2.mem[184][3] ),
    .A2(_01778_),
    .B(_01749_),
    .ZN(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06310_ (.A1(_01810_),
    .A2(_01811_),
    .A3(_01812_),
    .A4(_01813_),
    .ZN(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06311_ (.A1(\u2.mem[155][3] ),
    .A2(_01659_),
    .ZN(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06312_ (.A1(\u2.mem[174][3] ),
    .A2(_01656_),
    .B1(_01666_),
    .B2(\u2.mem[150][3] ),
    .C1(_01660_),
    .C2(\u2.mem[181][3] ),
    .ZN(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06313_ (.A1(\u2.mem[189][3] ),
    .A2(_01650_),
    .B1(_01652_),
    .B2(\u2.mem[176][3] ),
    .ZN(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06314_ (.A1(\u2.mem[172][3] ),
    .A2(_01654_),
    .B1(_01664_),
    .B2(\u2.mem[180][3] ),
    .ZN(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06315_ (.A1(_01815_),
    .A2(_01816_),
    .A3(_01817_),
    .A4(_01818_),
    .ZN(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06316_ (.A1(\u2.mem[177][3] ),
    .A2(_01734_),
    .B1(_01646_),
    .B2(\u2.mem[165][3] ),
    .C1(\u2.mem[163][3] ),
    .C2(_01642_),
    .ZN(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06317_ (.A1(\u2.mem[158][3] ),
    .A2(_01728_),
    .B1(_01729_),
    .B2(\u2.mem[151][3] ),
    .C1(_01731_),
    .C2(\u2.mem[193][3] ),
    .ZN(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06318_ (.A1(\u2.mem[145][3] ),
    .A2(_01640_),
    .B1(_01732_),
    .B2(\u2.mem[168][3] ),
    .ZN(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06319_ (.A1(\u2.mem[175][3] ),
    .A2(_01602_),
    .B1(_01631_),
    .B2(\u2.mem[188][3] ),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06320_ (.A1(\u2.mem[187][3] ),
    .A2(_01632_),
    .B1(_01635_),
    .B2(\u2.mem[192][3] ),
    .ZN(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06321_ (.A1(\u2.mem[159][3] ),
    .A2(_01604_),
    .B1(_01595_),
    .B2(\u2.mem[149][3] ),
    .ZN(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06322_ (.A1(_01823_),
    .A2(_01824_),
    .A3(_01825_),
    .ZN(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06323_ (.A1(\u2.mem[166][3] ),
    .A2(_01753_),
    .B1(_01754_),
    .B2(\u2.mem[161][3] ),
    .C(_01826_),
    .ZN(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06324_ (.A1(_01820_),
    .A2(_01821_),
    .A3(_01822_),
    .A4(_01827_),
    .ZN(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06325_ (.A1(\u2.mem[144][3] ),
    .A2(_01671_),
    .B1(_01673_),
    .B2(\u2.mem[182][3] ),
    .ZN(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06326_ (.A1(\u2.mem[190][3] ),
    .A2(_01702_),
    .B1(_01704_),
    .B2(\u2.mem[194][3] ),
    .ZN(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06327_ (.A1(\u2.mem[153][3] ),
    .A2(_01707_),
    .B1(_01709_),
    .B2(\u2.mem[160][3] ),
    .ZN(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06328_ (.A1(\u2.mem[152][3] ),
    .A2(_01712_),
    .B1(_01714_),
    .B2(\u2.mem[148][3] ),
    .ZN(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06329_ (.A1(_01830_),
    .A2(_01831_),
    .A3(_01832_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06330_ (.A1(\u2.mem[154][3] ),
    .A2(_01698_),
    .B1(_01700_),
    .B2(\u2.mem[162][3] ),
    .C(_01833_),
    .ZN(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06331_ (.A1(\u2.mem[173][3] ),
    .A2(_01720_),
    .B1(_01722_),
    .B2(\u2.mem[185][3] ),
    .ZN(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06332_ (.A1(\u2.mem[170][3] ),
    .A2(_01687_),
    .B1(_01689_),
    .B2(\u2.mem[156][3] ),
    .ZN(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06333_ (.A1(\u2.mem[191][3] ),
    .A2(_01682_),
    .B1(_01684_),
    .B2(\u2.mem[179][3] ),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06334_ (.A1(\u2.mem[146][3] ),
    .A2(_01692_),
    .B1(_01694_),
    .B2(\u2.mem[186][3] ),
    .ZN(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06335_ (.A1(_01836_),
    .A2(_01837_),
    .A3(_01838_),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06336_ (.A1(\u2.mem[147][3] ),
    .A2(_01676_),
    .B1(_01680_),
    .B2(\u2.mem[169][3] ),
    .C(_01839_),
    .ZN(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06337_ (.A1(_01829_),
    .A2(_01834_),
    .A3(_01835_),
    .A4(_01840_),
    .ZN(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06338_ (.A1(_01814_),
    .A2(_01819_),
    .A3(_01828_),
    .A4(_01841_),
    .ZN(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06339_ (.A1(_01809_),
    .A2(_01555_),
    .B(_01842_),
    .ZN(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06340_ (.I(\u2.mem[0][4] ),
    .ZN(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06341_ (.I(_01843_),
    .Z(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06342_ (.A1(\u2.mem[189][4] ),
    .A2(_01650_),
    .B1(_01663_),
    .B2(\u2.mem[180][4] ),
    .C1(_01652_),
    .C2(\u2.mem[176][4] ),
    .ZN(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06343_ (.A1(\u2.mem[174][4] ),
    .A2(_01657_),
    .B1(_01659_),
    .B2(\u2.mem[155][4] ),
    .C1(_01661_),
    .C2(\u2.mem[181][4] ),
    .ZN(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06344_ (.A1(\u2.mem[172][4] ),
    .A2(_01654_),
    .B1(_01667_),
    .B2(\u2.mem[150][4] ),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06345_ (.A1(_01845_),
    .A2(_01846_),
    .A3(_01847_),
    .ZN(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06346_ (.A1(\u2.mem[178][4] ),
    .A2(_01772_),
    .B1(_01773_),
    .B2(\u2.mem[164][4] ),
    .ZN(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06347_ (.A1(\u2.mem[167][4] ),
    .A2(_01775_),
    .B1(_01776_),
    .B2(\u2.mem[183][4] ),
    .ZN(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06348_ (.A1(\u2.mem[171][4] ),
    .A2(_01611_),
    .B1(_01770_),
    .B2(\u2.mem[157][4] ),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06349_ (.A1(\u2.mem[184][4] ),
    .A2(_01778_),
    .B(_01749_),
    .ZN(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06350_ (.A1(_01849_),
    .A2(_01850_),
    .A3(_01851_),
    .A4(_01852_),
    .ZN(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06351_ (.A1(\u2.mem[145][4] ),
    .A2(_01639_),
    .B1(_01643_),
    .B2(\u2.mem[163][4] ),
    .C1(\u2.mem[165][4] ),
    .C2(_01645_),
    .ZN(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06352_ (.A1(\u2.mem[158][4] ),
    .A2(_01728_),
    .B1(_01729_),
    .B2(\u2.mem[151][4] ),
    .C1(_01732_),
    .C2(\u2.mem[168][4] ),
    .ZN(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06353_ (.A1(\u2.mem[193][4] ),
    .A2(_01731_),
    .B1(_01734_),
    .B2(\u2.mem[177][4] ),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06354_ (.A1(\u2.mem[187][4] ),
    .A2(_01633_),
    .B1(_01636_),
    .B2(\u2.mem[192][4] ),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06355_ (.A1(\u2.mem[175][4] ),
    .A2(_01601_),
    .B1(_01630_),
    .B2(\u2.mem[188][4] ),
    .ZN(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06356_ (.A1(\u2.mem[159][4] ),
    .A2(_01603_),
    .B1(_01594_),
    .B2(\u2.mem[149][4] ),
    .ZN(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06357_ (.A1(_01857_),
    .A2(_01858_),
    .A3(_01859_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06358_ (.A1(\u2.mem[166][4] ),
    .A2(_01753_),
    .B1(_01754_),
    .B2(\u2.mem[161][4] ),
    .C(_01860_),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06359_ (.A1(_01854_),
    .A2(_01855_),
    .A3(_01856_),
    .A4(_01861_),
    .ZN(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06360_ (.A1(\u2.mem[190][4] ),
    .A2(_01703_),
    .B1(_01705_),
    .B2(\u2.mem[194][4] ),
    .ZN(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06361_ (.A1(\u2.mem[153][4] ),
    .A2(_01708_),
    .B1(_01710_),
    .B2(\u2.mem[160][4] ),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06362_ (.A1(\u2.mem[152][4] ),
    .A2(_01713_),
    .B1(_01715_),
    .B2(\u2.mem[148][4] ),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06363_ (.A1(_01863_),
    .A2(_01864_),
    .A3(_01865_),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06364_ (.A1(\u2.mem[154][4] ),
    .A2(_01699_),
    .B1(_01701_),
    .B2(\u2.mem[162][4] ),
    .C(_01866_),
    .ZN(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06365_ (.A1(\u2.mem[144][4] ),
    .A2(_01670_),
    .B1(_01672_),
    .B2(\u2.mem[182][4] ),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06366_ (.A1(\u2.mem[173][4] ),
    .A2(_01719_),
    .B1(_01721_),
    .B2(\u2.mem[185][4] ),
    .ZN(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06367_ (.A1(\u2.mem[170][4] ),
    .A2(_01686_),
    .B1(_01688_),
    .B2(\u2.mem[156][4] ),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06368_ (.A1(\u2.mem[191][4] ),
    .A2(_01681_),
    .B1(_01683_),
    .B2(\u2.mem[179][4] ),
    .ZN(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06369_ (.A1(\u2.mem[146][4] ),
    .A2(_01691_),
    .B1(_01693_),
    .B2(\u2.mem[186][4] ),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06370_ (.A1(_01870_),
    .A2(_01871_),
    .A3(_01872_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06371_ (.A1(\u2.mem[147][4] ),
    .A2(_01675_),
    .B1(_01679_),
    .B2(\u2.mem[169][4] ),
    .C(_01873_),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06372_ (.A1(_01867_),
    .A2(_01868_),
    .A3(_01869_),
    .A4(_01874_),
    .ZN(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06373_ (.A1(_01848_),
    .A2(_01853_),
    .A3(_01862_),
    .A4(_01875_),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06374_ (.A1(_01844_),
    .A2(_01555_),
    .B(_01876_),
    .ZN(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06375_ (.I(\u2.mem[0][5] ),
    .ZN(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06376_ (.I(_01877_),
    .Z(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06377_ (.A1(\u2.mem[189][5] ),
    .A2(_01650_),
    .B1(_01652_),
    .B2(\u2.mem[176][5] ),
    .C1(\u2.mem[172][5] ),
    .C2(_01653_),
    .ZN(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06378_ (.A1(\u2.mem[174][5] ),
    .A2(_01657_),
    .B1(_01659_),
    .B2(\u2.mem[155][5] ),
    .C1(_01661_),
    .C2(\u2.mem[181][5] ),
    .ZN(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06379_ (.A1(\u2.mem[180][5] ),
    .A2(_01664_),
    .B1(_01667_),
    .B2(\u2.mem[150][5] ),
    .ZN(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06380_ (.A1(_01879_),
    .A2(_01880_),
    .A3(_01881_),
    .ZN(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06381_ (.A1(\u2.mem[178][5] ),
    .A2(_01772_),
    .B1(_01773_),
    .B2(\u2.mem[164][5] ),
    .ZN(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06382_ (.A1(\u2.mem[167][5] ),
    .A2(_01775_),
    .B1(_01776_),
    .B2(\u2.mem[183][5] ),
    .ZN(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06383_ (.A1(\u2.mem[171][5] ),
    .A2(_01610_),
    .B1(_01770_),
    .B2(\u2.mem[157][5] ),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06384_ (.A1(\u2.mem[184][5] ),
    .A2(_01778_),
    .B(_01749_),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06385_ (.A1(_01883_),
    .A2(_01884_),
    .A3(_01885_),
    .A4(_01886_),
    .ZN(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06386_ (.A1(\u2.mem[177][5] ),
    .A2(_01583_),
    .B1(_01646_),
    .B2(\u2.mem[165][5] ),
    .C1(\u2.mem[163][5] ),
    .C2(_01642_),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06387_ (.A1(\u2.mem[158][5] ),
    .A2(_01728_),
    .B1(_01729_),
    .B2(\u2.mem[151][5] ),
    .C1(_01577_),
    .C2(\u2.mem[193][5] ),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06388_ (.A1(\u2.mem[145][5] ),
    .A2(_01640_),
    .B1(_01732_),
    .B2(\u2.mem[168][5] ),
    .ZN(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06389_ (.A1(\u2.mem[187][5] ),
    .A2(_01632_),
    .B1(_01635_),
    .B2(\u2.mem[192][5] ),
    .ZN(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06390_ (.A1(\u2.mem[175][5] ),
    .A2(_01601_),
    .B1(_01630_),
    .B2(\u2.mem[188][5] ),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06391_ (.A1(\u2.mem[159][5] ),
    .A2(_01603_),
    .B1(_01594_),
    .B2(\u2.mem[149][5] ),
    .ZN(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06392_ (.A1(_01891_),
    .A2(_01892_),
    .A3(_01893_),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06393_ (.A1(\u2.mem[166][5] ),
    .A2(_01592_),
    .B1(_01597_),
    .B2(\u2.mem[161][5] ),
    .C(_01894_),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06394_ (.A1(_01888_),
    .A2(_01889_),
    .A3(_01890_),
    .A4(_01895_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06395_ (.A1(\u2.mem[190][5] ),
    .A2(_01702_),
    .B1(_01704_),
    .B2(\u2.mem[194][5] ),
    .ZN(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06396_ (.A1(\u2.mem[153][5] ),
    .A2(_01707_),
    .B1(_01709_),
    .B2(\u2.mem[160][5] ),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06397_ (.A1(\u2.mem[152][5] ),
    .A2(_01712_),
    .B1(_01714_),
    .B2(\u2.mem[148][5] ),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06398_ (.A1(_01897_),
    .A2(_01898_),
    .A3(_01899_),
    .ZN(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06399_ (.A1(\u2.mem[154][5] ),
    .A2(_01699_),
    .B1(_01701_),
    .B2(\u2.mem[162][5] ),
    .C(_01900_),
    .ZN(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06400_ (.A1(\u2.mem[144][5] ),
    .A2(_01670_),
    .B1(_01672_),
    .B2(\u2.mem[182][5] ),
    .ZN(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06401_ (.A1(\u2.mem[173][5] ),
    .A2(_01719_),
    .B1(_01721_),
    .B2(\u2.mem[185][5] ),
    .ZN(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06402_ (.A1(\u2.mem[170][5] ),
    .A2(_01686_),
    .B1(_01688_),
    .B2(\u2.mem[156][5] ),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06403_ (.A1(\u2.mem[191][5] ),
    .A2(_01681_),
    .B1(_01683_),
    .B2(\u2.mem[179][5] ),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06404_ (.A1(\u2.mem[146][5] ),
    .A2(_01691_),
    .B1(_01693_),
    .B2(\u2.mem[186][5] ),
    .ZN(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06405_ (.A1(_01904_),
    .A2(_01905_),
    .A3(_01906_),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06406_ (.A1(\u2.mem[147][5] ),
    .A2(_01675_),
    .B1(_01679_),
    .B2(\u2.mem[169][5] ),
    .C(_01907_),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06407_ (.A1(_01901_),
    .A2(_01902_),
    .A3(_01903_),
    .A4(_01908_),
    .ZN(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06408_ (.A1(_01882_),
    .A2(_01887_),
    .A3(_01896_),
    .A4(_01909_),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06409_ (.A1(_01878_),
    .A2(_01554_),
    .B(_01910_),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06410_ (.I0(\u2.select_mem_row[5] ),
    .I1(\u2.select_mem_col[5] ),
    .S(_01510_),
    .Z(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06411_ (.I0(\u2.select_mem_row[4] ),
    .I1(\u2.select_mem_col[4] ),
    .S(_01502_),
    .Z(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06412_ (.A1(_01911_),
    .A2(_01912_),
    .Z(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06413_ (.I(_01913_),
    .Z(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06414_ (.I(_01914_),
    .Z(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06415_ (.I(_01912_),
    .Z(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06416_ (.I(_01916_),
    .Z(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06417_ (.A1(_01911_),
    .A2(_01916_),
    .ZN(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06418_ (.I(_01918_),
    .Z(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06419_ (.I(_01913_),
    .Z(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06420_ (.A1(\u2.mem[193][0] ),
    .A2(_01917_),
    .B1(_01919_),
    .B2(\u2.mem[192][0] ),
    .C(_01920_),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06421_ (.I(_01911_),
    .ZN(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06422_ (.A1(_01922_),
    .A2(_01916_),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06423_ (.I(_01923_),
    .Z(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06424_ (.A1(\u2.mem[194][0] ),
    .A2(_01924_),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06425_ (.A1(_01545_),
    .A2(_01915_),
    .B1(_01921_),
    .B2(_01925_),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06426_ (.A1(\u2.mem[194][1] ),
    .A2(_01924_),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06427_ (.I(_01916_),
    .Z(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06428_ (.I(_01927_),
    .Z(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06429_ (.I(_01918_),
    .Z(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06430_ (.A1(\u2.mem[193][1] ),
    .A2(_01928_),
    .B1(_01929_),
    .B2(\u2.mem[192][1] ),
    .C(_01914_),
    .ZN(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06431_ (.A1(_01727_),
    .A2(_01915_),
    .B1(_01926_),
    .B2(_01930_),
    .ZN(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06432_ (.I(_01919_),
    .Z(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06433_ (.A1(\u2.mem[192][2] ),
    .A2(_01931_),
    .ZN(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06434_ (.I(_01923_),
    .Z(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06435_ (.I(_01920_),
    .Z(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06436_ (.A1(\u2.mem[193][2] ),
    .A2(_01928_),
    .B1(_01933_),
    .B2(\u2.mem[194][2] ),
    .C(_01934_),
    .ZN(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06437_ (.A1(_01769_),
    .A2(_01915_),
    .B1(_01932_),
    .B2(_01935_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06438_ (.A1(\u2.mem[192][3] ),
    .A2(_01931_),
    .ZN(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06439_ (.A1(\u2.mem[193][3] ),
    .A2(_01928_),
    .B1(_01933_),
    .B2(\u2.mem[194][3] ),
    .C(_01934_),
    .ZN(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06440_ (.A1(_01809_),
    .A2(_01915_),
    .B1(_01936_),
    .B2(_01937_),
    .ZN(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06441_ (.I(_01914_),
    .Z(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06442_ (.A1(\u2.mem[194][4] ),
    .A2(_01924_),
    .ZN(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06443_ (.A1(\u2.mem[193][4] ),
    .A2(_01928_),
    .B1(_01929_),
    .B2(\u2.mem[192][4] ),
    .C(_01934_),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06444_ (.A1(_01844_),
    .A2(_01938_),
    .B1(_01939_),
    .B2(_01940_),
    .ZN(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06445_ (.A1(\u2.mem[192][5] ),
    .A2(_01931_),
    .ZN(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06446_ (.I(_01927_),
    .Z(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06447_ (.I(_01923_),
    .Z(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06448_ (.A1(\u2.mem[193][5] ),
    .A2(_01942_),
    .B1(_01943_),
    .B2(\u2.mem[194][5] ),
    .C(_01934_),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06449_ (.A1(_01878_),
    .A2(_01938_),
    .B1(_01941_),
    .B2(_01944_),
    .ZN(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06450_ (.I(\u2.mem[0][6] ),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06451_ (.I(_01923_),
    .Z(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06452_ (.A1(\u2.mem[194][6] ),
    .A2(_01946_),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06453_ (.I(_01918_),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06454_ (.I(_01913_),
    .Z(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06455_ (.A1(\u2.mem[193][6] ),
    .A2(_01942_),
    .B1(_01948_),
    .B2(\u2.mem[192][6] ),
    .C(_01949_),
    .ZN(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06456_ (.A1(_01945_),
    .A2(_01938_),
    .B1(_01947_),
    .B2(_01950_),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06457_ (.I(\u2.mem[0][7] ),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06458_ (.A1(\u2.mem[194][7] ),
    .A2(_01946_),
    .ZN(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06459_ (.A1(\u2.mem[193][7] ),
    .A2(_01942_),
    .B1(_01948_),
    .B2(\u2.mem[192][7] ),
    .C(_01949_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06460_ (.A1(_01951_),
    .A2(_01938_),
    .B1(_01952_),
    .B2(_01953_),
    .ZN(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06461_ (.I(\u2.mem[0][8] ),
    .ZN(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06462_ (.I(_01914_),
    .Z(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06463_ (.A1(\u2.mem[192][8] ),
    .A2(_01931_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06464_ (.A1(\u2.mem[193][8] ),
    .A2(_01942_),
    .B1(_01943_),
    .B2(\u2.mem[194][8] ),
    .C(_01949_),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06465_ (.A1(_01954_),
    .A2(_01955_),
    .B1(_01956_),
    .B2(_01957_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06466_ (.I(\u2.mem[0][9] ),
    .ZN(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06467_ (.A1(\u2.mem[192][9] ),
    .A2(_01929_),
    .ZN(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06468_ (.I(_01927_),
    .Z(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06469_ (.A1(\u2.mem[193][9] ),
    .A2(_01960_),
    .B1(_01943_),
    .B2(\u2.mem[194][9] ),
    .C(_01949_),
    .ZN(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06470_ (.A1(_01958_),
    .A2(_01955_),
    .B1(_01959_),
    .B2(_01961_),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06471_ (.I(\u2.mem[0][10] ),
    .ZN(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06472_ (.A1(\u2.mem[194][10] ),
    .A2(_01946_),
    .ZN(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06473_ (.I(_01913_),
    .Z(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06474_ (.A1(\u2.mem[193][10] ),
    .A2(_01960_),
    .B1(_01948_),
    .B2(\u2.mem[192][10] ),
    .C(_01964_),
    .ZN(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06475_ (.A1(_01962_),
    .A2(_01955_),
    .B1(_01963_),
    .B2(_01965_),
    .ZN(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06476_ (.I(\u2.mem[0][11] ),
    .ZN(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06477_ (.A1(\u2.mem[194][11] ),
    .A2(_01946_),
    .ZN(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06478_ (.A1(\u2.mem[193][11] ),
    .A2(_01960_),
    .B1(_01948_),
    .B2(\u2.mem[192][11] ),
    .C(_01964_),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06479_ (.A1(_01966_),
    .A2(_01955_),
    .B1(_01967_),
    .B2(_01968_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06480_ (.I(\u2.mem[0][12] ),
    .ZN(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06481_ (.I(_01920_),
    .Z(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06482_ (.A1(\u2.mem[192][12] ),
    .A2(_01929_),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06483_ (.A1(\u2.mem[193][12] ),
    .A2(_01960_),
    .B1(_01943_),
    .B2(\u2.mem[194][12] ),
    .C(_01964_),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06484_ (.A1(_01969_),
    .A2(_01970_),
    .B1(_01971_),
    .B2(_01972_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06485_ (.I(\u2.mem[0][13] ),
    .ZN(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06486_ (.A1(\u2.mem[194][13] ),
    .A2(_01933_),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06487_ (.A1(\u2.mem[193][13] ),
    .A2(_01917_),
    .B1(_01919_),
    .B2(\u2.mem[192][13] ),
    .C(_01964_),
    .ZN(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06488_ (.A1(_01973_),
    .A2(_01970_),
    .B1(_01974_),
    .B2(_01975_),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06489_ (.I(\u2.mem[0][14] ),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06490_ (.A1(\u2.mem[194][14] ),
    .A2(_01933_),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06491_ (.A1(\u2.mem[193][14] ),
    .A2(_01917_),
    .B1(_01919_),
    .B2(\u2.mem[192][14] ),
    .C(_01920_),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06492_ (.A1(_01976_),
    .A2(_01970_),
    .B1(_01977_),
    .B2(_01978_),
    .ZN(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06493_ (.I(\u2.mem[194][15] ),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06494_ (.I(\u2.mem[0][15] ),
    .ZN(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06495_ (.I(\u2.mem[192][15] ),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06496_ (.A1(_01981_),
    .A2(_01927_),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06497_ (.A1(\u2.mem[193][15] ),
    .A2(_01917_),
    .B(_01982_),
    .C(_01911_),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06498_ (.A1(_01979_),
    .A2(_01924_),
    .B1(_01970_),
    .B2(_01980_),
    .C(_01983_),
    .ZN(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06499_ (.I(\row_select_trans[0].data_sync ),
    .Z(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06500_ (.I(_01984_),
    .Z(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06501_ (.I(\row_select_trans[1].data_sync ),
    .Z(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06502_ (.A1(_01985_),
    .A2(_01986_),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06503_ (.I(\row_select_trans[2].data_sync ),
    .Z(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06504_ (.I(\row_select_trans[3].data_sync ),
    .Z(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06505_ (.A1(_01988_),
    .A2(_01989_),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06506_ (.I(_01990_),
    .Z(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06507_ (.A1(\row_select_trans[5].data_sync ),
    .A2(\row_select_trans[4].data_sync ),
    .ZN(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06508_ (.A1(_01987_),
    .A2(_01991_),
    .B(_01992_),
    .ZN(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06509_ (.I(_01993_),
    .Z(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06510_ (.I(_01994_),
    .Z(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06511_ (.I(_01995_),
    .Z(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06512_ (.I(\row_select_trans[4].data_sync ),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06513_ (.A1(\row_select_trans[5].data_sync ),
    .A2(_01997_),
    .ZN(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06514_ (.I(_01998_),
    .Z(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06515_ (.I(_01999_),
    .Z(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06516_ (.A1(_01985_),
    .A2(_01986_),
    .ZN(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06517_ (.A1(_01991_),
    .A2(_02001_),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06518_ (.A1(_02000_),
    .A2(_02002_),
    .ZN(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06519_ (.I(_02003_),
    .Z(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06520_ (.I(\row_select_trans[5].data_sync ),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06521_ (.A1(_02005_),
    .A2(\row_select_trans[4].data_sync ),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06522_ (.I(_02006_),
    .Z(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06523_ (.I(_01988_),
    .ZN(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06524_ (.I(_02008_),
    .Z(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06525_ (.I(\row_select_trans[3].data_sync ),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06526_ (.A1(_02009_),
    .A2(_02010_),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06527_ (.A1(_02011_),
    .A2(_02001_),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06528_ (.A1(_02007_),
    .A2(_02012_),
    .ZN(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06529_ (.I(_02013_),
    .Z(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06530_ (.I(_01998_),
    .Z(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06531_ (.I(_01984_),
    .ZN(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06532_ (.A1(_02016_),
    .A2(_01986_),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06533_ (.A1(_02017_),
    .A2(_02011_),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06534_ (.A1(_02015_),
    .A2(_02018_),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06535_ (.I(_02019_),
    .Z(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06536_ (.A1(\u2.mem[176][0] ),
    .A2(_02004_),
    .B1(_02014_),
    .B2(\u2.mem[172][0] ),
    .C1(_02020_),
    .C2(\u2.mem[189][0] ),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06537_ (.A1(_02005_),
    .A2(_01997_),
    .ZN(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06538_ (.I(_02022_),
    .Z(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06539_ (.I(\row_select_trans[1].data_sync ),
    .ZN(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06540_ (.I(_02024_),
    .Z(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06541_ (.A1(_02016_),
    .A2(_02025_),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06542_ (.A1(_01988_),
    .A2(_02010_),
    .ZN(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06543_ (.A1(_02026_),
    .A2(_02027_),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06544_ (.A1(_02023_),
    .A2(_02028_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06545_ (.I(_02029_),
    .Z(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06546_ (.I(_02006_),
    .Z(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06547_ (.A1(_01985_),
    .A2(_02025_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06548_ (.A1(_02032_),
    .A2(_02011_),
    .ZN(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06549_ (.A1(_02031_),
    .A2(_02033_),
    .ZN(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06550_ (.I(_02034_),
    .Z(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06551_ (.A1(_02009_),
    .A2(_01989_),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06552_ (.A1(_02017_),
    .A2(_02036_),
    .ZN(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06553_ (.A1(_02015_),
    .A2(_02037_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06554_ (.I(_02038_),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06555_ (.A1(\u2.mem[155][0] ),
    .A2(_02030_),
    .B1(_02035_),
    .B2(\u2.mem[174][0] ),
    .C1(\u2.mem[181][0] ),
    .C2(_02039_),
    .ZN(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06556_ (.A1(_02036_),
    .A2(_02001_),
    .ZN(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06557_ (.A1(_02041_),
    .A2(_02000_),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06558_ (.I(_02042_),
    .Z(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06559_ (.I(_02022_),
    .Z(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06560_ (.I(_02044_),
    .Z(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06561_ (.A1(_02032_),
    .A2(_02036_),
    .ZN(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06562_ (.A1(_02045_),
    .A2(_02046_),
    .ZN(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06563_ (.A1(\u2.mem[180][0] ),
    .A2(_02043_),
    .B1(_02047_),
    .B2(\u2.mem[150][0] ),
    .ZN(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06564_ (.A1(_02021_),
    .A2(_02040_),
    .A3(_02048_),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06565_ (.A1(_02031_),
    .A2(_02041_),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06566_ (.I(_02050_),
    .Z(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06567_ (.A1(_01990_),
    .A2(_02032_),
    .ZN(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06568_ (.I(_01998_),
    .Z(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06569_ (.A1(_02052_),
    .A2(_02053_),
    .ZN(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06570_ (.I(_02054_),
    .Z(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06571_ (.A1(\u2.mem[164][0] ),
    .A2(_02051_),
    .B1(_02055_),
    .B2(\u2.mem[178][0] ),
    .ZN(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06572_ (.I(_02006_),
    .Z(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06573_ (.A1(_02026_),
    .A2(_02036_),
    .ZN(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06574_ (.A1(_02057_),
    .A2(_02058_),
    .ZN(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06575_ (.I(_02059_),
    .Z(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06576_ (.A1(_02058_),
    .A2(_02053_),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06577_ (.I(_02061_),
    .Z(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06578_ (.A1(\u2.mem[167][0] ),
    .A2(_02060_),
    .B1(_02062_),
    .B2(\u2.mem[183][0] ),
    .ZN(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06579_ (.I(_02057_),
    .Z(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06580_ (.A1(_02064_),
    .A2(_02028_),
    .ZN(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06581_ (.I(_02065_),
    .Z(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06582_ (.A1(_02045_),
    .A2(_02018_),
    .ZN(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06583_ (.I(_02067_),
    .Z(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06584_ (.A1(\u2.mem[171][0] ),
    .A2(_02066_),
    .B1(_02068_),
    .B2(\u2.mem[157][0] ),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06585_ (.A1(_02027_),
    .A2(_02001_),
    .ZN(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06586_ (.A1(_02015_),
    .A2(_02070_),
    .ZN(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06587_ (.I(_02071_),
    .Z(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06588_ (.A1(\u2.mem[184][0] ),
    .A2(_02072_),
    .B(_01994_),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06589_ (.A1(_02056_),
    .A2(_02063_),
    .A3(_02069_),
    .A4(_02073_),
    .ZN(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06590_ (.A1(_02007_),
    .A2(_02037_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06591_ (.I(_02075_),
    .Z(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06592_ (.A1(_02026_),
    .A2(_01991_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06593_ (.A1(_02031_),
    .A2(_02077_),
    .ZN(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06594_ (.I(_02078_),
    .Z(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06595_ (.A1(_01991_),
    .A2(_02017_),
    .ZN(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06596_ (.A1(_02044_),
    .A2(_02080_),
    .ZN(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06597_ (.I(_02081_),
    .Z(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06598_ (.A1(\u2.mem[165][0] ),
    .A2(_02076_),
    .B1(_02079_),
    .B2(\u2.mem[163][0] ),
    .C1(\u2.mem[145][0] ),
    .C2(_02082_),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06599_ (.A1(_02023_),
    .A2(_02058_),
    .ZN(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06600_ (.I(_02084_),
    .Z(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06601_ (.A1(_02023_),
    .A2(_02033_),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06602_ (.I(_02086_),
    .Z(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06603_ (.A1(_01992_),
    .A2(_02080_),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06604_ (.I(_02088_),
    .Z(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06605_ (.A1(\u2.mem[151][0] ),
    .A2(_02085_),
    .B1(_02087_),
    .B2(\u2.mem[158][0] ),
    .C1(\u2.mem[193][0] ),
    .C2(_02089_),
    .ZN(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06606_ (.A1(_02080_),
    .A2(_02015_),
    .ZN(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06607_ (.I(_02091_),
    .Z(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06608_ (.A1(_02031_),
    .A2(_02070_),
    .ZN(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06609_ (.I(_02093_),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06610_ (.A1(\u2.mem[177][0] ),
    .A2(_02092_),
    .B1(_02094_),
    .B2(\u2.mem[168][0] ),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06611_ (.A1(_02064_),
    .A2(_02046_),
    .ZN(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06612_ (.I(_02096_),
    .Z(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06613_ (.A1(_02007_),
    .A2(_02080_),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06614_ (.I(_02098_),
    .Z(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06615_ (.A1(_02028_),
    .A2(_02053_),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06616_ (.A1(_01992_),
    .A2(_02002_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06617_ (.A1(\u2.mem[187][0] ),
    .A2(_02100_),
    .B1(_02101_),
    .B2(\u2.mem[192][0] ),
    .ZN(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06618_ (.A1(_02053_),
    .A2(_02012_),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06619_ (.A1(_02026_),
    .A2(_02011_),
    .ZN(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06620_ (.A1(_02057_),
    .A2(_02104_),
    .ZN(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06621_ (.A1(\u2.mem[188][0] ),
    .A2(_02103_),
    .B1(_02105_),
    .B2(\u2.mem[175][0] ),
    .ZN(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06622_ (.A1(_02044_),
    .A2(_02104_),
    .ZN(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06623_ (.I(_02022_),
    .Z(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06624_ (.A1(_02108_),
    .A2(_02037_),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06625_ (.A1(\u2.mem[159][0] ),
    .A2(_02107_),
    .B1(_02109_),
    .B2(\u2.mem[149][0] ),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06626_ (.A1(_02102_),
    .A2(_02106_),
    .A3(_02110_),
    .ZN(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06627_ (.A1(\u2.mem[166][0] ),
    .A2(_02097_),
    .B1(_02099_),
    .B2(\u2.mem[161][0] ),
    .C(_02111_),
    .ZN(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06628_ (.A1(_02083_),
    .A2(_02090_),
    .A3(_02095_),
    .A4(_02112_),
    .ZN(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06629_ (.A1(_02045_),
    .A2(_02002_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06630_ (.I(_02114_),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06631_ (.A1(_02000_),
    .A2(_02046_),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06632_ (.I(_02116_),
    .Z(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06633_ (.A1(\u2.mem[144][0] ),
    .A2(_02115_),
    .B1(_02117_),
    .B2(\u2.mem[182][0] ),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06634_ (.A1(_02027_),
    .A2(_02017_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06635_ (.A1(_02119_),
    .A2(_02000_),
    .ZN(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06636_ (.I(_02120_),
    .Z(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06637_ (.A1(_02064_),
    .A2(_02018_),
    .ZN(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06638_ (.I(_02122_),
    .Z(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06639_ (.A1(\u2.mem[185][0] ),
    .A2(_02121_),
    .B1(_02123_),
    .B2(\u2.mem[173][0] ),
    .ZN(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06640_ (.A1(_02027_),
    .A2(_02032_),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06641_ (.A1(_02045_),
    .A2(_02125_),
    .ZN(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06642_ (.A1(_02007_),
    .A2(_02052_),
    .ZN(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06643_ (.A1(_02108_),
    .A2(_02041_),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06644_ (.I(_02128_),
    .Z(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06645_ (.A1(_02108_),
    .A2(_02070_),
    .ZN(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06646_ (.I(_02130_),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06647_ (.A1(\u2.mem[148][0] ),
    .A2(_02129_),
    .B1(_02131_),
    .B2(\u2.mem[152][0] ),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06648_ (.A1(_01992_),
    .A2(_02052_),
    .ZN(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06649_ (.A1(_01999_),
    .A2(_02033_),
    .ZN(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06650_ (.A1(\u2.mem[194][0] ),
    .A2(_02133_),
    .B1(_02134_),
    .B2(\u2.mem[190][0] ),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06651_ (.A1(_02119_),
    .A2(_02044_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06652_ (.A1(_02006_),
    .A2(_02002_),
    .ZN(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06653_ (.A1(\u2.mem[153][0] ),
    .A2(_02136_),
    .B1(_02137_),
    .B2(\u2.mem[160][0] ),
    .ZN(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06654_ (.A1(_02132_),
    .A2(_02135_),
    .A3(_02138_),
    .ZN(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06655_ (.A1(\u2.mem[154][0] ),
    .A2(_02126_),
    .B1(_02127_),
    .B2(\u2.mem[162][0] ),
    .C(_02139_),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06656_ (.A1(_02064_),
    .A2(_02119_),
    .ZN(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06657_ (.I(_02141_),
    .Z(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06658_ (.A1(_02023_),
    .A2(_02077_),
    .ZN(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06659_ (.I(_02143_),
    .Z(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06660_ (.A1(_02057_),
    .A2(_02125_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06661_ (.I(_02145_),
    .Z(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06662_ (.A1(_02022_),
    .A2(_02012_),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06663_ (.I(_02147_),
    .Z(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06664_ (.A1(\u2.mem[170][0] ),
    .A2(_02146_),
    .B1(_02148_),
    .B2(\u2.mem[156][0] ),
    .ZN(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06665_ (.A1(_01998_),
    .A2(_02077_),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06666_ (.I(_02150_),
    .Z(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06667_ (.A1(_02104_),
    .A2(_01999_),
    .ZN(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06668_ (.I(_02152_),
    .Z(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06669_ (.A1(\u2.mem[179][0] ),
    .A2(_02151_),
    .B1(_02153_),
    .B2(\u2.mem[191][0] ),
    .ZN(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06670_ (.A1(_02108_),
    .A2(_02052_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06671_ (.I(_02155_),
    .Z(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06672_ (.A1(_02125_),
    .A2(_01999_),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06673_ (.I(_02157_),
    .Z(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06674_ (.A1(\u2.mem[146][0] ),
    .A2(_02156_),
    .B1(_02158_),
    .B2(\u2.mem[186][0] ),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06675_ (.A1(_02149_),
    .A2(_02154_),
    .A3(_02159_),
    .ZN(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06676_ (.A1(\u2.mem[169][0] ),
    .A2(_02142_),
    .B1(_02144_),
    .B2(\u2.mem[147][0] ),
    .C(_02160_),
    .ZN(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06677_ (.A1(_02118_),
    .A2(_02124_),
    .A3(_02140_),
    .A4(_02161_),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06678_ (.A1(_02049_),
    .A2(_02074_),
    .A3(_02113_),
    .A4(_02162_),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06679_ (.A1(_01545_),
    .A2(_01996_),
    .B(_02163_),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06680_ (.A1(\u2.mem[169][1] ),
    .A2(_02142_),
    .B1(_02144_),
    .B2(\u2.mem[147][1] ),
    .ZN(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06681_ (.A1(\u2.mem[144][1] ),
    .A2(_02115_),
    .B1(_02117_),
    .B2(\u2.mem[182][1] ),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06682_ (.A1(\u2.mem[185][1] ),
    .A2(_02121_),
    .B1(_02123_),
    .B2(\u2.mem[173][1] ),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06683_ (.A1(\u2.mem[170][1] ),
    .A2(_02146_),
    .B1(_02148_),
    .B2(\u2.mem[156][1] ),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06684_ (.A1(\u2.mem[179][1] ),
    .A2(_02151_),
    .B1(_02153_),
    .B2(\u2.mem[191][1] ),
    .ZN(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06685_ (.A1(_02167_),
    .A2(_02168_),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06686_ (.A1(\u2.mem[146][1] ),
    .A2(_02156_),
    .B1(_02158_),
    .B2(\u2.mem[186][1] ),
    .C(_02169_),
    .ZN(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06687_ (.A1(_02164_),
    .A2(_02165_),
    .A3(_02166_),
    .A4(_02170_),
    .Z(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06688_ (.A1(\u2.mem[151][1] ),
    .A2(_02085_),
    .B1(_02087_),
    .B2(\u2.mem[158][1] ),
    .C1(\u2.mem[193][1] ),
    .C2(_02089_),
    .ZN(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06689_ (.A1(\u2.mem[145][1] ),
    .A2(_02082_),
    .B1(_02094_),
    .B2(\u2.mem[168][1] ),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06690_ (.I(_02107_),
    .Z(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06691_ (.A1(\u2.mem[166][1] ),
    .A2(_02096_),
    .B1(_02098_),
    .B2(\u2.mem[161][1] ),
    .C1(\u2.mem[159][1] ),
    .C2(_02174_),
    .ZN(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06692_ (.I(_02109_),
    .Z(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06693_ (.I(_02105_),
    .Z(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06694_ (.A1(\u2.mem[149][1] ),
    .A2(_02176_),
    .B1(_02177_),
    .B2(\u2.mem[175][1] ),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06695_ (.A1(_02172_),
    .A2(_02173_),
    .A3(_02175_),
    .A4(_02178_),
    .ZN(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06696_ (.A1(\u2.mem[164][1] ),
    .A2(_02050_),
    .B1(_02054_),
    .B2(\u2.mem[178][1] ),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06697_ (.A1(\u2.mem[167][1] ),
    .A2(_02059_),
    .B1(_02061_),
    .B2(\u2.mem[183][1] ),
    .ZN(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06698_ (.A1(\u2.mem[184][1] ),
    .A2(_02071_),
    .B(_01993_),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06699_ (.A1(_02180_),
    .A2(_02181_),
    .A3(_02182_),
    .ZN(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06700_ (.A1(\u2.mem[171][1] ),
    .A2(_02065_),
    .B1(_02067_),
    .B2(\u2.mem[157][1] ),
    .C(_02183_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06701_ (.I(_02103_),
    .Z(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06702_ (.I(_02100_),
    .Z(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06703_ (.I(_02101_),
    .Z(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06704_ (.A1(\u2.mem[188][1] ),
    .A2(_02185_),
    .B1(_02186_),
    .B2(\u2.mem[187][1] ),
    .C1(_02187_),
    .C2(\u2.mem[192][1] ),
    .ZN(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06705_ (.A1(\u2.mem[165][1] ),
    .A2(_02076_),
    .B1(_02079_),
    .B2(\u2.mem[163][1] ),
    .C1(_02092_),
    .C2(\u2.mem[177][1] ),
    .ZN(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06706_ (.A1(_02184_),
    .A2(_02188_),
    .A3(_02189_),
    .ZN(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06707_ (.A1(\u2.mem[155][1] ),
    .A2(_02030_),
    .B1(_02035_),
    .B2(\u2.mem[174][1] ),
    .C1(\u2.mem[181][1] ),
    .C2(_02039_),
    .ZN(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06708_ (.I(_02047_),
    .Z(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06709_ (.A1(\u2.mem[180][1] ),
    .A2(_02043_),
    .B1(_02192_),
    .B2(\u2.mem[150][1] ),
    .ZN(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06710_ (.A1(_02191_),
    .A2(_02193_),
    .ZN(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06711_ (.A1(\u2.mem[154][1] ),
    .A2(_02126_),
    .B1(_02129_),
    .B2(\u2.mem[148][1] ),
    .C1(_02127_),
    .C2(\u2.mem[162][1] ),
    .ZN(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06712_ (.I(_02136_),
    .Z(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06713_ (.A1(\u2.mem[153][1] ),
    .A2(_02196_),
    .B1(_02131_),
    .B2(\u2.mem[152][1] ),
    .ZN(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06714_ (.I(_02133_),
    .Z(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06715_ (.I(_02134_),
    .Z(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06716_ (.I(_02137_),
    .Z(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06717_ (.A1(\u2.mem[194][1] ),
    .A2(_02198_),
    .B1(_02199_),
    .B2(\u2.mem[190][1] ),
    .C1(_02200_),
    .C2(\u2.mem[160][1] ),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _06718_ (.A1(\u2.mem[176][1] ),
    .A2(_02003_),
    .B1(_02013_),
    .B2(\u2.mem[172][1] ),
    .C1(_02019_),
    .C2(\u2.mem[189][1] ),
    .ZN(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06719_ (.A1(_02195_),
    .A2(_02197_),
    .A3(_02201_),
    .A4(_02202_),
    .ZN(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06720_ (.A1(_02179_),
    .A2(_02190_),
    .A3(_02194_),
    .A4(_02203_),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06721_ (.A1(_01727_),
    .A2(_01995_),
    .B1(_02171_),
    .B2(_02204_),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06722_ (.A1(\u2.mem[164][2] ),
    .A2(_02051_),
    .B1(_02055_),
    .B2(\u2.mem[178][2] ),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06723_ (.A1(\u2.mem[167][2] ),
    .A2(_02060_),
    .B1(_02062_),
    .B2(\u2.mem[183][2] ),
    .ZN(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06724_ (.A1(\u2.mem[171][2] ),
    .A2(_02066_),
    .B1(_02068_),
    .B2(\u2.mem[157][2] ),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06725_ (.A1(\u2.mem[184][2] ),
    .A2(_02072_),
    .B(_01995_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06726_ (.A1(_02205_),
    .A2(_02206_),
    .A3(_02207_),
    .A4(_02208_),
    .ZN(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06727_ (.A1(\u2.mem[150][2] ),
    .A2(_02192_),
    .ZN(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06728_ (.A1(\u2.mem[155][2] ),
    .A2(_02030_),
    .B1(_02035_),
    .B2(\u2.mem[174][2] ),
    .C1(\u2.mem[181][2] ),
    .C2(_02039_),
    .ZN(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06729_ (.A1(\u2.mem[176][2] ),
    .A2(_02004_),
    .B1(_02020_),
    .B2(\u2.mem[189][2] ),
    .ZN(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06730_ (.A1(\u2.mem[180][2] ),
    .A2(_02043_),
    .B1(_02014_),
    .B2(\u2.mem[172][2] ),
    .ZN(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06731_ (.A1(_02210_),
    .A2(_02211_),
    .A3(_02212_),
    .A4(_02213_),
    .ZN(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06732_ (.A1(\u2.mem[187][2] ),
    .A2(_02186_),
    .B1(_02187_),
    .B2(\u2.mem[192][2] ),
    .ZN(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06733_ (.A1(\u2.mem[188][2] ),
    .A2(_02185_),
    .B1(_02177_),
    .B2(\u2.mem[175][2] ),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06734_ (.A1(\u2.mem[159][2] ),
    .A2(_02174_),
    .B1(_02176_),
    .B2(\u2.mem[149][2] ),
    .ZN(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06735_ (.A1(_02215_),
    .A2(_02216_),
    .A3(_02217_),
    .ZN(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06736_ (.A1(\u2.mem[166][2] ),
    .A2(_02097_),
    .B1(_02099_),
    .B2(\u2.mem[161][2] ),
    .C(_02218_),
    .ZN(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06737_ (.A1(\u2.mem[165][2] ),
    .A2(_02076_),
    .B1(_02079_),
    .B2(\u2.mem[163][2] ),
    .C1(\u2.mem[145][2] ),
    .C2(_02081_),
    .ZN(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06738_ (.A1(\u2.mem[151][2] ),
    .A2(_02085_),
    .B1(_02087_),
    .B2(\u2.mem[158][2] ),
    .C1(\u2.mem[168][2] ),
    .C2(_02094_),
    .ZN(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06739_ (.A1(\u2.mem[177][2] ),
    .A2(_02092_),
    .B1(_02089_),
    .B2(\u2.mem[193][2] ),
    .ZN(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06740_ (.A1(_02219_),
    .A2(_02220_),
    .A3(_02221_),
    .A4(_02222_),
    .ZN(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06741_ (.A1(\u2.mem[144][2] ),
    .A2(_02115_),
    .B1(_02117_),
    .B2(\u2.mem[182][2] ),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06742_ (.I(_02126_),
    .Z(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06743_ (.I(_02127_),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06744_ (.A1(\u2.mem[194][2] ),
    .A2(_02198_),
    .B1(_02199_),
    .B2(\u2.mem[190][2] ),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06745_ (.A1(\u2.mem[153][2] ),
    .A2(_02196_),
    .B1(_02200_),
    .B2(\u2.mem[160][2] ),
    .ZN(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06746_ (.A1(\u2.mem[148][2] ),
    .A2(_02128_),
    .B1(_02130_),
    .B2(\u2.mem[152][2] ),
    .ZN(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06747_ (.A1(_02227_),
    .A2(_02228_),
    .A3(_02229_),
    .ZN(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06748_ (.A1(\u2.mem[154][2] ),
    .A2(_02225_),
    .B1(_02226_),
    .B2(\u2.mem[162][2] ),
    .C(_02230_),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06749_ (.A1(\u2.mem[185][2] ),
    .A2(_02121_),
    .B1(_02123_),
    .B2(\u2.mem[173][2] ),
    .ZN(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06750_ (.A1(\u2.mem[170][2] ),
    .A2(_02145_),
    .B1(_02147_),
    .B2(\u2.mem[156][2] ),
    .ZN(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06751_ (.A1(\u2.mem[179][2] ),
    .A2(_02150_),
    .B1(_02152_),
    .B2(\u2.mem[191][2] ),
    .ZN(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06752_ (.A1(\u2.mem[146][2] ),
    .A2(_02155_),
    .B1(_02157_),
    .B2(\u2.mem[186][2] ),
    .ZN(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06753_ (.A1(_02233_),
    .A2(_02234_),
    .A3(_02235_),
    .ZN(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06754_ (.A1(\u2.mem[169][2] ),
    .A2(_02141_),
    .B1(_02143_),
    .B2(\u2.mem[147][2] ),
    .C(_02236_),
    .ZN(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06755_ (.A1(_02224_),
    .A2(_02231_),
    .A3(_02232_),
    .A4(_02237_),
    .ZN(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06756_ (.A1(_02209_),
    .A2(_02214_),
    .A3(_02223_),
    .A4(_02238_),
    .ZN(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06757_ (.A1(_01769_),
    .A2(_01996_),
    .B(_02239_),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06758_ (.A1(\u2.mem[159][3] ),
    .A2(_02174_),
    .B1(_02176_),
    .B2(\u2.mem[149][3] ),
    .ZN(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06759_ (.A1(\u2.mem[187][3] ),
    .A2(_02186_),
    .B1(_02187_),
    .B2(\u2.mem[192][3] ),
    .ZN(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06760_ (.A1(\u2.mem[188][3] ),
    .A2(_02185_),
    .B1(_02177_),
    .B2(\u2.mem[175][3] ),
    .ZN(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06761_ (.A1(_02240_),
    .A2(_02241_),
    .A3(_02242_),
    .ZN(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06762_ (.A1(\u2.mem[166][3] ),
    .A2(_02097_),
    .B1(_02099_),
    .B2(\u2.mem[161][3] ),
    .C(_02243_),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06763_ (.A1(\u2.mem[154][3] ),
    .A2(_02225_),
    .B1(_02226_),
    .B2(\u2.mem[162][3] ),
    .ZN(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06764_ (.A1(\u2.mem[194][3] ),
    .A2(_02198_),
    .B1(_02199_),
    .B2(\u2.mem[190][3] ),
    .ZN(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06765_ (.A1(\u2.mem[153][3] ),
    .A2(_02196_),
    .B1(_02200_),
    .B2(\u2.mem[160][3] ),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06766_ (.A1(_02246_),
    .A2(_02247_),
    .ZN(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06767_ (.A1(\u2.mem[148][3] ),
    .A2(_02129_),
    .B1(_02131_),
    .B2(\u2.mem[152][3] ),
    .C(_02248_),
    .ZN(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06768_ (.A1(\u2.mem[169][3] ),
    .A2(_02142_),
    .B1(_02144_),
    .B2(\u2.mem[147][3] ),
    .C1(_02158_),
    .C2(\u2.mem[186][3] ),
    .ZN(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06769_ (.A1(\u2.mem[164][3] ),
    .A2(_02051_),
    .B1(_02055_),
    .B2(\u2.mem[178][3] ),
    .ZN(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06770_ (.A1(\u2.mem[167][3] ),
    .A2(_02060_),
    .B1(_02062_),
    .B2(\u2.mem[183][3] ),
    .ZN(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06771_ (.A1(\u2.mem[171][3] ),
    .A2(_02065_),
    .B1(_02067_),
    .B2(\u2.mem[157][3] ),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06772_ (.A1(\u2.mem[184][3] ),
    .A2(_02072_),
    .B(_01994_),
    .ZN(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06773_ (.A1(_02251_),
    .A2(_02252_),
    .A3(_02253_),
    .A4(_02254_),
    .ZN(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06774_ (.A1(\u2.mem[168][3] ),
    .A2(_02093_),
    .ZN(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06775_ (.A1(\u2.mem[151][3] ),
    .A2(_02084_),
    .B1(_02086_),
    .B2(\u2.mem[158][3] ),
    .C1(\u2.mem[193][3] ),
    .C2(_02088_),
    .ZN(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06776_ (.A1(\u2.mem[165][3] ),
    .A2(_02075_),
    .B1(_02078_),
    .B2(\u2.mem[163][3] ),
    .ZN(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06777_ (.A1(\u2.mem[145][3] ),
    .A2(_02081_),
    .B1(_02091_),
    .B2(\u2.mem[177][3] ),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06778_ (.A1(_02256_),
    .A2(_02257_),
    .A3(_02258_),
    .A4(_02259_),
    .ZN(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06779_ (.A1(\u2.mem[180][3] ),
    .A2(_02042_),
    .B1(_02013_),
    .B2(\u2.mem[172][3] ),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06780_ (.A1(\u2.mem[155][3] ),
    .A2(_02029_),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06781_ (.A1(\u2.mem[150][3] ),
    .A2(_02047_),
    .B1(_02034_),
    .B2(\u2.mem[174][3] ),
    .C1(\u2.mem[181][3] ),
    .C2(_02038_),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06782_ (.A1(\u2.mem[176][3] ),
    .A2(_02003_),
    .B1(_02019_),
    .B2(\u2.mem[189][3] ),
    .ZN(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06783_ (.A1(_02261_),
    .A2(_02262_),
    .A3(_02263_),
    .A4(_02264_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06784_ (.A1(\u2.mem[170][3] ),
    .A2(_02146_),
    .B1(_02148_),
    .B2(\u2.mem[156][3] ),
    .ZN(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06785_ (.A1(\u2.mem[179][3] ),
    .A2(_02151_),
    .B1(_02153_),
    .B2(\u2.mem[191][3] ),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06786_ (.A1(\u2.mem[185][3] ),
    .A2(_02120_),
    .B1(_02116_),
    .B2(\u2.mem[182][3] ),
    .C1(\u2.mem[144][3] ),
    .C2(_02114_),
    .ZN(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06787_ (.A1(\u2.mem[146][3] ),
    .A2(_02156_),
    .B1(_02122_),
    .B2(\u2.mem[173][3] ),
    .ZN(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06788_ (.A1(_02266_),
    .A2(_02267_),
    .A3(_02268_),
    .A4(_02269_),
    .ZN(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06789_ (.A1(_02255_),
    .A2(_02260_),
    .A3(_02265_),
    .A4(_02270_),
    .ZN(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06790_ (.A1(_02245_),
    .A2(_02249_),
    .A3(_02250_),
    .A4(_02271_),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06791_ (.A1(_01809_),
    .A2(_01995_),
    .B1(_02244_),
    .B2(_02272_),
    .ZN(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06792_ (.A1(\u2.mem[151][4] ),
    .A2(_02084_),
    .B1(_02086_),
    .B2(\u2.mem[158][4] ),
    .C1(\u2.mem[168][4] ),
    .C2(_02093_),
    .ZN(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06793_ (.A1(\u2.mem[177][4] ),
    .A2(_02091_),
    .B1(_02088_),
    .B2(\u2.mem[193][4] ),
    .ZN(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06794_ (.A1(\u2.mem[166][4] ),
    .A2(_02096_),
    .B1(_02098_),
    .B2(\u2.mem[161][4] ),
    .C1(\u2.mem[159][4] ),
    .C2(_02174_),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06795_ (.A1(\u2.mem[149][4] ),
    .A2(_02176_),
    .B1(_02177_),
    .B2(\u2.mem[175][4] ),
    .ZN(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06796_ (.A1(_02273_),
    .A2(_02274_),
    .A3(_02275_),
    .A4(_02276_),
    .Z(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06797_ (.A1(\u2.mem[164][4] ),
    .A2(_02050_),
    .B1(_02054_),
    .B2(\u2.mem[178][4] ),
    .ZN(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06798_ (.A1(\u2.mem[167][4] ),
    .A2(_02059_),
    .B1(_02061_),
    .B2(\u2.mem[183][4] ),
    .ZN(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06799_ (.A1(\u2.mem[184][4] ),
    .A2(_02071_),
    .B(_01993_),
    .ZN(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06800_ (.A1(_02278_),
    .A2(_02279_),
    .A3(_02280_),
    .ZN(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06801_ (.A1(\u2.mem[171][4] ),
    .A2(_02066_),
    .B1(_02068_),
    .B2(\u2.mem[157][4] ),
    .C(_02281_),
    .ZN(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06802_ (.A1(\u2.mem[188][4] ),
    .A2(_02185_),
    .B1(_02186_),
    .B2(\u2.mem[187][4] ),
    .C1(_02187_),
    .C2(\u2.mem[192][4] ),
    .ZN(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06803_ (.A1(\u2.mem[165][4] ),
    .A2(_02076_),
    .B1(_02079_),
    .B2(\u2.mem[163][4] ),
    .C1(\u2.mem[145][4] ),
    .C2(_02082_),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06804_ (.A1(_02277_),
    .A2(_02282_),
    .A3(_02283_),
    .A4(_02284_),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06805_ (.A1(\u2.mem[176][4] ),
    .A2(_02004_),
    .B1(_02020_),
    .B2(\u2.mem[189][4] ),
    .ZN(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06806_ (.A1(\u2.mem[180][4] ),
    .A2(_02043_),
    .B1(_02014_),
    .B2(\u2.mem[172][4] ),
    .ZN(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06807_ (.A1(\u2.mem[174][4] ),
    .A2(_02035_),
    .B1(_02039_),
    .B2(\u2.mem[181][4] ),
    .ZN(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06808_ (.A1(\u2.mem[155][4] ),
    .A2(_02030_),
    .B1(_02192_),
    .B2(\u2.mem[150][4] ),
    .ZN(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06809_ (.A1(_02286_),
    .A2(_02287_),
    .A3(_02288_),
    .A4(_02289_),
    .ZN(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06810_ (.A1(\u2.mem[146][4] ),
    .A2(_02156_),
    .B1(_02158_),
    .B2(\u2.mem[186][4] ),
    .ZN(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06811_ (.A1(\u2.mem[170][4] ),
    .A2(_02146_),
    .B1(_02148_),
    .B2(\u2.mem[156][4] ),
    .ZN(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06812_ (.A1(\u2.mem[179][4] ),
    .A2(_02151_),
    .B1(_02153_),
    .B2(\u2.mem[191][4] ),
    .ZN(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06813_ (.A1(_02291_),
    .A2(_02292_),
    .A3(_02293_),
    .ZN(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06814_ (.A1(\u2.mem[169][4] ),
    .A2(_02142_),
    .B1(_02144_),
    .B2(\u2.mem[147][4] ),
    .C(_02294_),
    .ZN(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06815_ (.A1(\u2.mem[194][4] ),
    .A2(_02198_),
    .B1(_02199_),
    .B2(\u2.mem[190][4] ),
    .ZN(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06816_ (.A1(\u2.mem[153][4] ),
    .A2(_02196_),
    .B1(_02200_),
    .B2(\u2.mem[160][4] ),
    .ZN(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06817_ (.A1(\u2.mem[148][4] ),
    .A2(_02129_),
    .B1(_02131_),
    .B2(\u2.mem[152][4] ),
    .ZN(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06818_ (.A1(_02296_),
    .A2(_02297_),
    .A3(_02298_),
    .ZN(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06819_ (.A1(\u2.mem[154][4] ),
    .A2(_02225_),
    .B1(_02226_),
    .B2(\u2.mem[162][4] ),
    .C(_02299_),
    .ZN(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06820_ (.A1(\u2.mem[144][4] ),
    .A2(_02115_),
    .B1(_02117_),
    .B2(\u2.mem[182][4] ),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06821_ (.A1(\u2.mem[185][4] ),
    .A2(_02121_),
    .B1(_02123_),
    .B2(\u2.mem[173][4] ),
    .ZN(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06822_ (.A1(_02295_),
    .A2(_02300_),
    .A3(_02301_),
    .A4(_02302_),
    .ZN(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06823_ (.A1(_02285_),
    .A2(_02290_),
    .A3(_02303_),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06824_ (.A1(_01844_),
    .A2(_01996_),
    .B(_02304_),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06825_ (.A1(\u2.mem[171][5] ),
    .A2(_02066_),
    .B1(_02068_),
    .B2(\u2.mem[157][5] ),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06826_ (.A1(\u2.mem[164][5] ),
    .A2(_02051_),
    .B1(_02055_),
    .B2(\u2.mem[178][5] ),
    .ZN(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06827_ (.A1(\u2.mem[167][5] ),
    .A2(_02060_),
    .B1(_02062_),
    .B2(\u2.mem[183][5] ),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06828_ (.A1(\u2.mem[184][5] ),
    .A2(_02072_),
    .B(_01994_),
    .ZN(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06829_ (.A1(_02305_),
    .A2(_02306_),
    .A3(_02307_),
    .A4(_02308_),
    .ZN(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06830_ (.A1(\u2.mem[150][5] ),
    .A2(_02192_),
    .ZN(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06831_ (.A1(\u2.mem[155][5] ),
    .A2(_02029_),
    .B1(_02034_),
    .B2(\u2.mem[174][5] ),
    .C1(\u2.mem[181][5] ),
    .C2(_02038_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06832_ (.A1(\u2.mem[176][5] ),
    .A2(_02004_),
    .B1(_02020_),
    .B2(\u2.mem[189][5] ),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06833_ (.A1(\u2.mem[180][5] ),
    .A2(_02042_),
    .B1(_02014_),
    .B2(\u2.mem[172][5] ),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06834_ (.A1(_02310_),
    .A2(_02311_),
    .A3(_02312_),
    .A4(_02313_),
    .ZN(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06835_ (.A1(\u2.mem[187][5] ),
    .A2(_02100_),
    .B1(_02101_),
    .B2(\u2.mem[192][5] ),
    .ZN(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06836_ (.A1(\u2.mem[188][5] ),
    .A2(_02103_),
    .B1(_02105_),
    .B2(\u2.mem[175][5] ),
    .ZN(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06837_ (.A1(\u2.mem[159][5] ),
    .A2(_02107_),
    .B1(_02109_),
    .B2(\u2.mem[149][5] ),
    .ZN(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06838_ (.A1(_02315_),
    .A2(_02316_),
    .A3(_02317_),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06839_ (.A1(\u2.mem[166][5] ),
    .A2(_02097_),
    .B1(_02099_),
    .B2(\u2.mem[161][5] ),
    .C(_02318_),
    .ZN(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06840_ (.A1(\u2.mem[165][5] ),
    .A2(_02075_),
    .B1(_02078_),
    .B2(\u2.mem[163][5] ),
    .C1(_02092_),
    .C2(\u2.mem[177][5] ),
    .ZN(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06841_ (.A1(\u2.mem[151][5] ),
    .A2(_02085_),
    .B1(_02087_),
    .B2(\u2.mem[158][5] ),
    .C1(\u2.mem[193][5] ),
    .C2(_02089_),
    .ZN(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06842_ (.A1(\u2.mem[145][5] ),
    .A2(_02082_),
    .B1(_02094_),
    .B2(\u2.mem[168][5] ),
    .ZN(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06843_ (.A1(_02319_),
    .A2(_02320_),
    .A3(_02321_),
    .A4(_02322_),
    .ZN(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06844_ (.A1(\u2.mem[144][5] ),
    .A2(_02114_),
    .B1(_02116_),
    .B2(\u2.mem[182][5] ),
    .ZN(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06845_ (.A1(\u2.mem[194][5] ),
    .A2(_02133_),
    .B1(_02134_),
    .B2(\u2.mem[190][5] ),
    .ZN(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06846_ (.A1(\u2.mem[153][5] ),
    .A2(_02136_),
    .B1(_02137_),
    .B2(\u2.mem[160][5] ),
    .ZN(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06847_ (.A1(\u2.mem[148][5] ),
    .A2(_02128_),
    .B1(_02130_),
    .B2(\u2.mem[152][5] ),
    .ZN(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06848_ (.A1(_02325_),
    .A2(_02326_),
    .A3(_02327_),
    .ZN(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06849_ (.A1(\u2.mem[154][5] ),
    .A2(_02225_),
    .B1(_02226_),
    .B2(\u2.mem[162][5] ),
    .C(_02328_),
    .ZN(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06850_ (.A1(\u2.mem[185][5] ),
    .A2(_02120_),
    .B1(_02122_),
    .B2(\u2.mem[173][5] ),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06851_ (.A1(\u2.mem[170][5] ),
    .A2(_02145_),
    .B1(_02147_),
    .B2(\u2.mem[156][5] ),
    .ZN(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06852_ (.A1(\u2.mem[179][5] ),
    .A2(_02150_),
    .B1(_02152_),
    .B2(\u2.mem[191][5] ),
    .ZN(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06853_ (.A1(\u2.mem[146][5] ),
    .A2(_02155_),
    .B1(_02157_),
    .B2(\u2.mem[186][5] ),
    .ZN(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06854_ (.A1(_02331_),
    .A2(_02332_),
    .A3(_02333_),
    .ZN(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06855_ (.A1(\u2.mem[169][5] ),
    .A2(_02141_),
    .B1(_02143_),
    .B2(\u2.mem[147][5] ),
    .C(_02334_),
    .ZN(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06856_ (.A1(_02324_),
    .A2(_02329_),
    .A3(_02330_),
    .A4(_02335_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06857_ (.A1(_02309_),
    .A2(_02314_),
    .A3(_02323_),
    .A4(_02336_),
    .ZN(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06858_ (.A1(_01878_),
    .A2(_01996_),
    .B(_02337_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06859_ (.A1(_02009_),
    .A2(\row_select_trans[4].data_sync ),
    .Z(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06860_ (.A1(_02025_),
    .A2(_01989_),
    .ZN(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06861_ (.A1(\row_select_trans[0].data_sync ),
    .A2(\row_select_trans[2].data_sync ),
    .Z(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06862_ (.A1(\col_select_trans[5].data_sync ),
    .A2(_02025_),
    .ZN(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06863_ (.A1(\col_select_trans[5].data_sync ),
    .A2(_02024_),
    .B(_02016_),
    .C(\col_select_trans[4].data_sync ),
    .ZN(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06864_ (.A1(_01984_),
    .A2(_02008_),
    .B1(_02010_),
    .B2(\row_select_trans[1].data_sync ),
    .ZN(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06865_ (.A1(_02340_),
    .A2(_02341_),
    .A3(_02342_),
    .B(_02343_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06866_ (.A1(_02339_),
    .A2(_02344_),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06867_ (.A1(_02338_),
    .A2(_02345_),
    .Z(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06868_ (.I(_02346_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06869_ (.A1(_01579_),
    .A2(_01985_),
    .Z(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06870_ (.I(_02348_),
    .ZN(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06871_ (.A1(\col_select_trans[5].data_sync ),
    .A2(_01986_),
    .Z(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06872_ (.A1(_02349_),
    .A2(_02350_),
    .ZN(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06873_ (.I(_02340_),
    .Z(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06874_ (.A1(_01989_),
    .A2(\row_select_trans[5].data_sync ),
    .Z(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06875_ (.A1(\row_select_trans[1].data_sync ),
    .A2(_02010_),
    .ZN(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06876_ (.A1(_02339_),
    .A2(_02354_),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06877_ (.A1(_02352_),
    .A2(_02353_),
    .A3(_02355_),
    .ZN(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06878_ (.A1(_02347_),
    .A2(_02351_),
    .A3(_02356_),
    .Z(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06879_ (.I(_02357_),
    .Z(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06880_ (.I(_02358_),
    .Z(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06881_ (.I(_02359_),
    .Z(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06882_ (.I(_02360_),
    .Z(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06883_ (.A1(_02338_),
    .A2(_02345_),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06884_ (.I(_02362_),
    .Z(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06885_ (.I(_02363_),
    .Z(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06886_ (.A1(_01988_),
    .A2(_01997_),
    .ZN(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06887_ (.I(_02365_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06888_ (.A1(_02339_),
    .A2(_02338_),
    .A3(_02344_),
    .Z(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06889_ (.I(_02353_),
    .ZN(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06890_ (.A1(_02366_),
    .A2(_02367_),
    .A3(_02368_),
    .ZN(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06891_ (.I(_02369_),
    .Z(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06892_ (.I(_02370_),
    .Z(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06893_ (.A1(_02339_),
    .A2(_02338_),
    .A3(_02344_),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06894_ (.A1(_02365_),
    .A2(_02372_),
    .B(_02353_),
    .ZN(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06895_ (.I(_02373_),
    .Z(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _06896_ (.I(_02374_),
    .Z(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06897_ (.A1(_02341_),
    .A2(_02342_),
    .ZN(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06898_ (.A1(_02352_),
    .A2(_02376_),
    .Z(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06899_ (.I(_02377_),
    .Z(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06900_ (.A1(_01984_),
    .A2(_02009_),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _06901_ (.A1(_02352_),
    .A2(_02341_),
    .A3(_02342_),
    .B(_02379_),
    .ZN(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06902_ (.A1(_02355_),
    .A2(_02380_),
    .Z(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06903_ (.I(_02381_),
    .Z(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06904_ (.I(_02351_),
    .Z(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06905_ (.A1(_02378_),
    .A2(_02382_),
    .A3(_02383_),
    .ZN(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06906_ (.A1(_02364_),
    .A2(_02371_),
    .A3(_02375_),
    .A4(_02384_),
    .ZN(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06907_ (.I(_02385_),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06908_ (.A1(_02365_),
    .A2(_02372_),
    .A3(_02353_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _06909_ (.I(_02387_),
    .Z(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06910_ (.A1(_02366_),
    .A2(_02367_),
    .B(_02368_),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _06911_ (.I(_02389_),
    .Z(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06912_ (.I(_02381_),
    .Z(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06913_ (.A1(_02348_),
    .A2(_02350_),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06914_ (.A1(_02378_),
    .A2(_02391_),
    .A3(_02392_),
    .ZN(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06915_ (.I(_02363_),
    .Z(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06916_ (.A1(_02388_),
    .A2(_02390_),
    .B(_02393_),
    .C(_02394_),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06917_ (.I(_02395_),
    .Z(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06918_ (.A1(\u2.mem[32][0] ),
    .A2(_02386_),
    .B1(_02396_),
    .B2(\u2.mem[2][0] ),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06919_ (.I(_02363_),
    .Z(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06920_ (.I(_02370_),
    .Z(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _06921_ (.I(_02374_),
    .Z(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06922_ (.I(_02377_),
    .Z(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06923_ (.A1(_02355_),
    .A2(_02380_),
    .ZN(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06924_ (.I(_02402_),
    .Z(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06925_ (.A1(_02401_),
    .A2(_02403_),
    .A3(_02383_),
    .ZN(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06926_ (.A1(_02398_),
    .A2(_02399_),
    .A3(_02400_),
    .A4(_02404_),
    .ZN(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06927_ (.I(_02405_),
    .Z(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06928_ (.I(_02387_),
    .Z(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06929_ (.I(_02389_),
    .Z(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06930_ (.A1(_02352_),
    .A2(_02376_),
    .ZN(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06931_ (.I(_02409_),
    .Z(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06932_ (.A1(_02410_),
    .A2(_02403_),
    .A3(_02392_),
    .ZN(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06933_ (.I(_02346_),
    .Z(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06934_ (.I(_02412_),
    .Z(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06935_ (.A1(_02407_),
    .A2(_02408_),
    .B(_02411_),
    .C(_02413_),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06936_ (.I(_02414_),
    .Z(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06937_ (.A1(\u2.mem[40][0] ),
    .A2(_02406_),
    .B1(_02415_),
    .B2(\u2.mem[30][0] ),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06938_ (.I(_02387_),
    .Z(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06939_ (.I(_02417_),
    .Z(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06940_ (.I(_02389_),
    .Z(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06941_ (.I(_02419_),
    .Z(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06942_ (.I(_02402_),
    .Z(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06943_ (.A1(_01551_),
    .A2(_02016_),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06944_ (.A1(_02422_),
    .A2(_02350_),
    .Z(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06945_ (.A1(_02349_),
    .A2(_02423_),
    .Z(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06946_ (.A1(_02378_),
    .A2(_02421_),
    .A3(_02424_),
    .ZN(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06947_ (.I(_02412_),
    .Z(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06948_ (.A1(_02418_),
    .A2(_02420_),
    .B(_02425_),
    .C(_02426_),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06949_ (.I(_02427_),
    .Z(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06950_ (.I(_02362_),
    .Z(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06951_ (.I(_02369_),
    .Z(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06952_ (.I(_02430_),
    .Z(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06953_ (.I(_02373_),
    .Z(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06954_ (.I(_02432_),
    .Z(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06955_ (.A1(_02401_),
    .A2(_02391_),
    .A3(_02424_),
    .ZN(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06956_ (.A1(_02429_),
    .A2(_02431_),
    .A3(_02433_),
    .A4(_02434_),
    .ZN(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06957_ (.I(_02435_),
    .Z(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06958_ (.A1(\u2.mem[27][0] ),
    .A2(_02428_),
    .B1(_02436_),
    .B2(\u2.mem[35][0] ),
    .ZN(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06959_ (.I(_02370_),
    .Z(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _06960_ (.I(_02374_),
    .Z(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06961_ (.A1(_02348_),
    .A2(_02423_),
    .ZN(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06962_ (.I(_02409_),
    .Z(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06963_ (.A1(_02440_),
    .A2(_02441_),
    .A3(_02421_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06964_ (.A1(_02398_),
    .A2(_02438_),
    .A3(_02439_),
    .A4(_02442_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06965_ (.I(_02443_),
    .Z(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06966_ (.I(_02430_),
    .Z(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06967_ (.I(_02432_),
    .Z(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06968_ (.A1(_02429_),
    .A2(_02445_),
    .A3(_02446_),
    .A4(_02393_),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06969_ (.I(_02447_),
    .Z(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06970_ (.A1(\u2.mem[45][0] ),
    .A2(_02444_),
    .B1(_02448_),
    .B2(\u2.mem[34][0] ),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06971_ (.A1(_02397_),
    .A2(_02416_),
    .A3(_02437_),
    .A4(_02449_),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06972_ (.I(_02407_),
    .Z(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06973_ (.I(_02408_),
    .Z(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06974_ (.A1(_02441_),
    .A2(_02421_),
    .A3(_02424_),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06975_ (.I(_02362_),
    .Z(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06976_ (.I(_02454_),
    .Z(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06977_ (.A1(_02451_),
    .A2(_02452_),
    .B(_02453_),
    .C(_02455_),
    .ZN(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06978_ (.I(_02456_),
    .Z(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06979_ (.I(_02417_),
    .Z(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06980_ (.I(_02419_),
    .Z(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06981_ (.A1(_02458_),
    .A2(_02459_),
    .B(_02442_),
    .C(_02364_),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06982_ (.I(_02460_),
    .Z(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06983_ (.A1(\u2.mem[15][0] ),
    .A2(_02457_),
    .B1(_02461_),
    .B2(\u2.mem[13][0] ),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06984_ (.A1(_02440_),
    .A2(_02401_),
    .A3(_02382_),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06985_ (.A1(_02458_),
    .A2(_02459_),
    .B(_02463_),
    .C(_02398_),
    .ZN(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06986_ (.I(_02464_),
    .Z(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06987_ (.I(_02387_),
    .Z(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06988_ (.I(_02389_),
    .Z(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06989_ (.A1(_02410_),
    .A2(_02391_),
    .A3(_02424_),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06990_ (.I(_02362_),
    .Z(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06991_ (.A1(_02466_),
    .A2(_02467_),
    .B(_02468_),
    .C(_02469_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06992_ (.I(_02470_),
    .Z(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06993_ (.A1(\u2.mem[1][0] ),
    .A2(_02465_),
    .B1(_02471_),
    .B2(\u2.mem[7][0] ),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06994_ (.I(_02412_),
    .Z(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06995_ (.A1(_02388_),
    .A2(_02390_),
    .B(_02384_),
    .C(_02473_),
    .ZN(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06996_ (.I(_02474_),
    .Z(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06997_ (.A1(_02429_),
    .A2(_02445_),
    .A3(_02446_),
    .A4(_02463_),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06998_ (.I(_02476_),
    .Z(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06999_ (.A1(\u2.mem[16][0] ),
    .A2(_02475_),
    .B1(_02477_),
    .B2(\u2.mem[33][0] ),
    .ZN(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07000_ (.A1(_02451_),
    .A2(_02452_),
    .B(_02434_),
    .C(_02455_),
    .ZN(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07001_ (.I(_02479_),
    .Z(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07002_ (.A1(\u2.mem[3][0] ),
    .A2(_02480_),
    .B(_02359_),
    .ZN(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07003_ (.A1(_02462_),
    .A2(_02472_),
    .A3(_02478_),
    .A4(_02481_),
    .ZN(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07004_ (.I(_02412_),
    .Z(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07005_ (.A1(_02440_),
    .A2(_02441_),
    .A3(_02382_),
    .ZN(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07006_ (.A1(_02483_),
    .A2(_02438_),
    .A3(_02439_),
    .A4(_02484_),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07007_ (.I(_02485_),
    .Z(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07008_ (.I(_02346_),
    .Z(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07009_ (.A1(_02487_),
    .A2(_02445_),
    .A3(_02446_),
    .A4(_02404_),
    .ZN(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07010_ (.I(_02488_),
    .Z(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07011_ (.A1(\u2.mem[53][0] ),
    .A2(_02486_),
    .B1(_02489_),
    .B2(\u2.mem[56][0] ),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07012_ (.I(_02430_),
    .Z(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _07013_ (.I(_02432_),
    .Z(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07014_ (.A1(_02401_),
    .A2(_02403_),
    .A3(_02392_),
    .ZN(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07015_ (.A1(_02413_),
    .A2(_02491_),
    .A3(_02492_),
    .A4(_02493_),
    .ZN(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07016_ (.I(_02494_),
    .Z(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07017_ (.I(_02430_),
    .Z(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _07018_ (.I(_02432_),
    .Z(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07019_ (.A1(_02410_),
    .A2(_02391_),
    .A3(_02383_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07020_ (.A1(_02454_),
    .A2(_02496_),
    .A3(_02497_),
    .A4(_02498_),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07021_ (.I(_02499_),
    .Z(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07022_ (.A1(\u2.mem[58][0] ),
    .A2(_02495_),
    .B1(_02500_),
    .B2(\u2.mem[36][0] ),
    .ZN(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07023_ (.A1(_02483_),
    .A2(_02491_),
    .A3(_02492_),
    .A4(_02393_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07024_ (.I(_02502_),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07025_ (.A1(_02487_),
    .A2(_02496_),
    .A3(_02497_),
    .A4(_02434_),
    .ZN(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07026_ (.I(_02504_),
    .Z(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07027_ (.A1(\u2.mem[50][0] ),
    .A2(_02503_),
    .B1(_02505_),
    .B2(\u2.mem[51][0] ),
    .ZN(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07028_ (.A1(_02441_),
    .A2(_02382_),
    .A3(_02392_),
    .ZN(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07029_ (.A1(_02413_),
    .A2(_02491_),
    .A3(_02492_),
    .A4(_02507_),
    .ZN(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07030_ (.I(_02508_),
    .Z(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07031_ (.A1(_02487_),
    .A2(_02496_),
    .A3(_02497_),
    .A4(_02468_),
    .ZN(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07032_ (.I(_02510_),
    .Z(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07033_ (.A1(\u2.mem[54][0] ),
    .A2(_02509_),
    .B1(_02511_),
    .B2(\u2.mem[55][0] ),
    .ZN(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07034_ (.A1(_02490_),
    .A2(_02501_),
    .A3(_02506_),
    .A4(_02512_),
    .ZN(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07035_ (.A1(_02469_),
    .A2(_02431_),
    .A3(_02433_),
    .A4(_02425_),
    .ZN(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07036_ (.I(_02514_),
    .Z(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07037_ (.A1(_02407_),
    .A2(_02408_),
    .B(_02498_),
    .C(_02487_),
    .ZN(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07038_ (.I(_02516_),
    .Z(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07039_ (.A1(\u2.mem[43][0] ),
    .A2(_02515_),
    .B1(_02517_),
    .B2(\u2.mem[20][0] ),
    .ZN(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07040_ (.A1(_02410_),
    .A2(_02403_),
    .A3(_02383_),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07041_ (.A1(_02394_),
    .A2(_02438_),
    .A3(_02439_),
    .A4(_02519_),
    .ZN(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07042_ (.I(_02520_),
    .Z(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _07043_ (.A1(_02429_),
    .A2(_02445_),
    .A3(_02446_),
    .A4(_02493_),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07044_ (.I(_02522_),
    .Z(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07045_ (.A1(\u2.mem[44][0] ),
    .A2(_02521_),
    .B1(_02523_),
    .B2(\u2.mem[42][0] ),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07046_ (.A1(_02466_),
    .A2(_02467_),
    .B(_02411_),
    .C(_02394_),
    .ZN(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07047_ (.I(_02525_),
    .Z(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07048_ (.A1(_02407_),
    .A2(_02408_),
    .B(_02519_),
    .C(_02454_),
    .ZN(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07049_ (.I(_02527_),
    .Z(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07050_ (.A1(\u2.mem[14][0] ),
    .A2(_02526_),
    .B1(_02528_),
    .B2(\u2.mem[12][0] ),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07051_ (.A1(_02413_),
    .A2(_02431_),
    .A3(_02433_),
    .A4(_02463_),
    .ZN(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07052_ (.I(_02530_),
    .Z(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07053_ (.A1(_02454_),
    .A2(_02496_),
    .A3(_02497_),
    .A4(_02411_),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07054_ (.I(_02532_),
    .Z(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07055_ (.A1(\u2.mem[49][0] ),
    .A2(_02531_),
    .B1(_02533_),
    .B2(\u2.mem[46][0] ),
    .ZN(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07056_ (.A1(_02518_),
    .A2(_02524_),
    .A3(_02529_),
    .A4(_02534_),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07057_ (.A1(_02450_),
    .A2(_02482_),
    .A3(_02513_),
    .A4(_02535_),
    .ZN(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07058_ (.I(_02370_),
    .Z(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _07059_ (.I(_02374_),
    .Z(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07060_ (.A1(_02455_),
    .A2(_02537_),
    .A3(_02538_),
    .A4(_02484_),
    .ZN(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07061_ (.I(_02539_),
    .Z(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07062_ (.A1(_02426_),
    .A2(_02399_),
    .A3(_02400_),
    .A4(_02425_),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07063_ (.I(_02541_),
    .Z(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07064_ (.A1(\u2.mem[37][0] ),
    .A2(_02540_),
    .B1(_02542_),
    .B2(\u2.mem[59][0] ),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07065_ (.I(_02347_),
    .Z(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07066_ (.A1(_02544_),
    .A2(_02537_),
    .A3(_02538_),
    .A4(_02519_),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07067_ (.I(_02545_),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07068_ (.I(_02347_),
    .Z(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07069_ (.A1(_02547_),
    .A2(_02371_),
    .A3(_02375_),
    .A4(_02411_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07070_ (.I(_02548_),
    .Z(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07071_ (.A1(\u2.mem[60][0] ),
    .A2(_02546_),
    .B1(_02549_),
    .B2(\u2.mem[62][0] ),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07072_ (.I(_02347_),
    .Z(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07073_ (.A1(_02440_),
    .A2(_02378_),
    .A3(_02421_),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07074_ (.A1(_02551_),
    .A2(_02537_),
    .A3(_02538_),
    .A4(_02552_),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07075_ (.I(_02553_),
    .Z(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07076_ (.A1(_02398_),
    .A2(_02399_),
    .A3(_02400_),
    .A4(_02552_),
    .ZN(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07077_ (.I(_02555_),
    .Z(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07078_ (.A1(\u2.mem[57][0] ),
    .A2(_02554_),
    .B1(_02556_),
    .B2(\u2.mem[41][0] ),
    .ZN(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07079_ (.A1(_02551_),
    .A2(_02537_),
    .A3(_02538_),
    .A4(_02442_),
    .ZN(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07080_ (.I(_02558_),
    .Z(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07081_ (.A1(_02473_),
    .A2(_02399_),
    .A3(_02400_),
    .A4(_02453_),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07082_ (.I(_02560_),
    .Z(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07083_ (.A1(\u2.mem[61][0] ),
    .A2(_02559_),
    .B1(_02561_),
    .B2(\u2.mem[63][0] ),
    .ZN(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07084_ (.A1(_02543_),
    .A2(_02550_),
    .A3(_02557_),
    .A4(_02562_),
    .ZN(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07085_ (.A1(_02451_),
    .A2(_02452_),
    .B(_02442_),
    .C(_02544_),
    .ZN(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07086_ (.I(_02564_),
    .Z(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07087_ (.I(_02417_),
    .Z(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07088_ (.I(_02419_),
    .Z(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07089_ (.I(_02363_),
    .Z(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07090_ (.A1(_02566_),
    .A2(_02567_),
    .B(_02425_),
    .C(_02568_),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07091_ (.I(_02569_),
    .Z(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07092_ (.A1(\u2.mem[29][0] ),
    .A2(_02565_),
    .B1(_02570_),
    .B2(\u2.mem[11][0] ),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07093_ (.A1(_02451_),
    .A2(_02452_),
    .B(_02493_),
    .C(_02544_),
    .ZN(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07094_ (.I(_02572_),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07095_ (.A1(_02566_),
    .A2(_02567_),
    .B(_02493_),
    .C(_02568_),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07096_ (.I(_02574_),
    .Z(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07097_ (.A1(\u2.mem[26][0] ),
    .A2(_02573_),
    .B1(_02575_),
    .B2(\u2.mem[10][0] ),
    .ZN(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07098_ (.I(_02417_),
    .Z(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07099_ (.I(_02419_),
    .Z(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07100_ (.A1(_02577_),
    .A2(_02578_),
    .B(_02552_),
    .C(_02455_),
    .ZN(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07101_ (.I(_02579_),
    .Z(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07102_ (.A1(_02418_),
    .A2(_02420_),
    .B(_02552_),
    .C(_02426_),
    .ZN(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07103_ (.I(_02581_),
    .Z(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07104_ (.A1(\u2.mem[9][0] ),
    .A2(_02580_),
    .B1(_02582_),
    .B2(\u2.mem[25][0] ),
    .ZN(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07105_ (.A1(_02577_),
    .A2(_02578_),
    .B(_02519_),
    .C(_02551_),
    .ZN(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07106_ (.I(_02584_),
    .Z(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07107_ (.A1(_02388_),
    .A2(_02390_),
    .B(_02453_),
    .C(_02473_),
    .ZN(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07108_ (.I(_02586_),
    .Z(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07109_ (.A1(\u2.mem[28][0] ),
    .A2(_02585_),
    .B1(_02587_),
    .B2(\u2.mem[31][0] ),
    .ZN(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07110_ (.A1(_02571_),
    .A2(_02576_),
    .A3(_02583_),
    .A4(_02588_),
    .ZN(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07111_ (.A1(_02577_),
    .A2(_02578_),
    .B(_02463_),
    .C(_02544_),
    .ZN(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07112_ (.I(_02590_),
    .Z(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07113_ (.A1(_02418_),
    .A2(_02420_),
    .B(_02404_),
    .C(_02547_),
    .ZN(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07114_ (.I(_02592_),
    .Z(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07115_ (.A1(\u2.mem[17][0] ),
    .A2(_02591_),
    .B1(_02593_),
    .B2(\u2.mem[24][0] ),
    .ZN(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07116_ (.A1(_02577_),
    .A2(_02578_),
    .B(_02468_),
    .C(_02551_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07117_ (.I(_02595_),
    .Z(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07118_ (.A1(_02418_),
    .A2(_02420_),
    .B(_02507_),
    .C(_02426_),
    .ZN(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07119_ (.I(_02597_),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07120_ (.A1(\u2.mem[23][0] ),
    .A2(_02596_),
    .B1(_02598_),
    .B2(\u2.mem[22][0] ),
    .ZN(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07121_ (.A1(_02547_),
    .A2(_02371_),
    .A3(_02375_),
    .A4(_02498_),
    .ZN(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07122_ (.I(_02600_),
    .Z(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07123_ (.A1(_02388_),
    .A2(_02390_),
    .B(_02484_),
    .C(_02483_),
    .ZN(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07124_ (.I(_02602_),
    .Z(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07125_ (.A1(\u2.mem[52][0] ),
    .A2(_02601_),
    .B1(_02603_),
    .B2(\u2.mem[21][0] ),
    .ZN(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07126_ (.A1(_02566_),
    .A2(_02567_),
    .B(_02393_),
    .C(_02547_),
    .ZN(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07127_ (.I(_02605_),
    .Z(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07128_ (.A1(_02466_),
    .A2(_02467_),
    .B(_02434_),
    .C(_02483_),
    .ZN(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07129_ (.I(_02607_),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07130_ (.A1(\u2.mem[18][0] ),
    .A2(_02606_),
    .B1(_02608_),
    .B2(\u2.mem[19][0] ),
    .ZN(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07131_ (.A1(_02594_),
    .A2(_02599_),
    .A3(_02604_),
    .A4(_02609_),
    .ZN(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07132_ (.A1(_02566_),
    .A2(_02567_),
    .B(_02404_),
    .C(_02568_),
    .ZN(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07133_ (.I(_02611_),
    .Z(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07134_ (.A1(_02466_),
    .A2(_02467_),
    .B(_02498_),
    .C(_02394_),
    .ZN(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07135_ (.I(_02613_),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07136_ (.A1(\u2.mem[8][0] ),
    .A2(_02612_),
    .B1(_02614_),
    .B2(\u2.mem[4][0] ),
    .ZN(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07137_ (.A1(_02568_),
    .A2(_02371_),
    .A3(_02375_),
    .A4(_02468_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07138_ (.I(_02616_),
    .Z(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07139_ (.A1(_02473_),
    .A2(_02438_),
    .A3(_02439_),
    .A4(_02384_),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07140_ (.I(_02618_),
    .Z(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07141_ (.A1(\u2.mem[39][0] ),
    .A2(_02617_),
    .B1(_02619_),
    .B2(\u2.mem[48][0] ),
    .ZN(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07142_ (.A1(_02458_),
    .A2(_02459_),
    .B(_02507_),
    .C(_02364_),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07143_ (.I(_02621_),
    .Z(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07144_ (.A1(_02469_),
    .A2(_02491_),
    .A3(_02492_),
    .A4(_02453_),
    .ZN(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07145_ (.I(_02623_),
    .Z(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07146_ (.A1(\u2.mem[6][0] ),
    .A2(_02622_),
    .B1(_02624_),
    .B2(\u2.mem[47][0] ),
    .ZN(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07147_ (.A1(_02458_),
    .A2(_02459_),
    .B(_02484_),
    .C(_02364_),
    .ZN(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07148_ (.I(_02626_),
    .Z(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _07149_ (.A1(_02469_),
    .A2(_02431_),
    .A3(_02433_),
    .A4(_02507_),
    .ZN(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07150_ (.I(_02628_),
    .Z(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07151_ (.A1(\u2.mem[5][0] ),
    .A2(_02627_),
    .B1(_02629_),
    .B2(\u2.mem[38][0] ),
    .ZN(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07152_ (.A1(_02615_),
    .A2(_02620_),
    .A3(_02625_),
    .A4(_02630_),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07153_ (.A1(_02563_),
    .A2(_02589_),
    .A3(_02610_),
    .A4(_02631_),
    .ZN(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07154_ (.A1(_01544_),
    .A2(_02361_),
    .B1(_02536_),
    .B2(_02632_),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07155_ (.I(_02443_),
    .Z(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07156_ (.I(_02447_),
    .Z(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07157_ (.A1(\u2.mem[45][1] ),
    .A2(_02633_),
    .B1(_02634_),
    .B2(\u2.mem[34][1] ),
    .ZN(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07158_ (.A1(\u2.mem[32][1] ),
    .A2(_02386_),
    .B1(_02396_),
    .B2(\u2.mem[2][1] ),
    .ZN(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07159_ (.A1(\u2.mem[40][1] ),
    .A2(_02406_),
    .B1(_02415_),
    .B2(\u2.mem[30][1] ),
    .ZN(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07160_ (.A1(\u2.mem[27][1] ),
    .A2(_02428_),
    .B1(_02436_),
    .B2(\u2.mem[35][1] ),
    .ZN(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07161_ (.A1(_02635_),
    .A2(_02636_),
    .A3(_02637_),
    .A4(_02638_),
    .ZN(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07162_ (.A1(\u2.mem[15][1] ),
    .A2(_02457_),
    .B1(_02461_),
    .B2(\u2.mem[13][1] ),
    .ZN(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07163_ (.A1(\u2.mem[1][1] ),
    .A2(_02465_),
    .B1(_02471_),
    .B2(\u2.mem[7][1] ),
    .ZN(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07164_ (.A1(\u2.mem[16][1] ),
    .A2(_02475_),
    .B1(_02477_),
    .B2(\u2.mem[33][1] ),
    .ZN(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07165_ (.A1(\u2.mem[3][1] ),
    .A2(_02480_),
    .B(_02359_),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07166_ (.A1(_02640_),
    .A2(_02641_),
    .A3(_02642_),
    .A4(_02643_),
    .ZN(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07167_ (.I(_02502_),
    .Z(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07168_ (.I(_02504_),
    .Z(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07169_ (.A1(\u2.mem[50][1] ),
    .A2(_02645_),
    .B1(_02646_),
    .B2(\u2.mem[51][1] ),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07170_ (.I(_02508_),
    .Z(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07171_ (.I(_02510_),
    .Z(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07172_ (.A1(\u2.mem[54][1] ),
    .A2(_02648_),
    .B1(_02649_),
    .B2(\u2.mem[55][1] ),
    .ZN(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07173_ (.A1(\u2.mem[53][1] ),
    .A2(_02486_),
    .B1(_02489_),
    .B2(\u2.mem[56][1] ),
    .ZN(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07174_ (.A1(\u2.mem[58][1] ),
    .A2(_02495_),
    .B1(_02500_),
    .B2(\u2.mem[36][1] ),
    .ZN(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07175_ (.A1(_02647_),
    .A2(_02650_),
    .A3(_02651_),
    .A4(_02652_),
    .ZN(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07176_ (.I(_02520_),
    .Z(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07177_ (.I(_02522_),
    .Z(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07178_ (.A1(\u2.mem[44][1] ),
    .A2(_02654_),
    .B1(_02655_),
    .B2(\u2.mem[42][1] ),
    .ZN(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07179_ (.I(_02525_),
    .Z(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07180_ (.I(_02527_),
    .Z(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07181_ (.A1(\u2.mem[14][1] ),
    .A2(_02657_),
    .B1(_02658_),
    .B2(\u2.mem[12][1] ),
    .ZN(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07182_ (.I(_02530_),
    .Z(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07183_ (.I(_02532_),
    .Z(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07184_ (.A1(\u2.mem[49][1] ),
    .A2(_02660_),
    .B1(_02661_),
    .B2(\u2.mem[46][1] ),
    .ZN(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07185_ (.A1(\u2.mem[43][1] ),
    .A2(_02515_),
    .B1(_02517_),
    .B2(\u2.mem[20][1] ),
    .ZN(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07186_ (.A1(_02656_),
    .A2(_02659_),
    .A3(_02662_),
    .A4(_02663_),
    .ZN(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07187_ (.A1(_02639_),
    .A2(_02644_),
    .A3(_02653_),
    .A4(_02664_),
    .ZN(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07188_ (.I(_02558_),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07189_ (.I(_02560_),
    .Z(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07190_ (.A1(\u2.mem[61][1] ),
    .A2(_02666_),
    .B1(_02667_),
    .B2(\u2.mem[63][1] ),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07191_ (.A1(\u2.mem[60][1] ),
    .A2(_02546_),
    .B1(_02549_),
    .B2(\u2.mem[62][1] ),
    .ZN(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07192_ (.A1(\u2.mem[37][1] ),
    .A2(_02540_),
    .B1(_02542_),
    .B2(\u2.mem[59][1] ),
    .ZN(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07193_ (.A1(\u2.mem[57][1] ),
    .A2(_02554_),
    .B1(_02556_),
    .B2(\u2.mem[41][1] ),
    .ZN(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07194_ (.A1(_02668_),
    .A2(_02669_),
    .A3(_02670_),
    .A4(_02671_),
    .ZN(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07195_ (.I(_02572_),
    .Z(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07196_ (.I(_02574_),
    .Z(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07197_ (.A1(\u2.mem[26][1] ),
    .A2(_02673_),
    .B1(_02674_),
    .B2(\u2.mem[10][1] ),
    .ZN(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07198_ (.A1(\u2.mem[29][1] ),
    .A2(_02565_),
    .B1(_02570_),
    .B2(\u2.mem[11][1] ),
    .ZN(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07199_ (.A1(\u2.mem[9][1] ),
    .A2(_02580_),
    .B1(_02582_),
    .B2(\u2.mem[25][1] ),
    .ZN(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07200_ (.A1(\u2.mem[28][1] ),
    .A2(_02585_),
    .B1(_02587_),
    .B2(\u2.mem[31][1] ),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07201_ (.A1(_02675_),
    .A2(_02676_),
    .A3(_02677_),
    .A4(_02678_),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07202_ (.I(_02595_),
    .Z(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07203_ (.I(_02597_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07204_ (.A1(\u2.mem[23][1] ),
    .A2(_02680_),
    .B1(_02681_),
    .B2(\u2.mem[22][1] ),
    .ZN(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07205_ (.A1(\u2.mem[17][1] ),
    .A2(_02591_),
    .B1(_02593_),
    .B2(\u2.mem[24][1] ),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07206_ (.A1(\u2.mem[52][1] ),
    .A2(_02601_),
    .B1(_02603_),
    .B2(\u2.mem[21][1] ),
    .ZN(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07207_ (.A1(\u2.mem[18][1] ),
    .A2(_02606_),
    .B1(_02608_),
    .B2(\u2.mem[19][1] ),
    .ZN(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07208_ (.A1(_02682_),
    .A2(_02683_),
    .A3(_02684_),
    .A4(_02685_),
    .ZN(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07209_ (.I(_02626_),
    .Z(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07210_ (.I(_02628_),
    .Z(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07211_ (.A1(\u2.mem[5][1] ),
    .A2(_02687_),
    .B1(_02688_),
    .B2(\u2.mem[38][1] ),
    .ZN(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07212_ (.A1(\u2.mem[39][1] ),
    .A2(_02617_),
    .B1(_02619_),
    .B2(\u2.mem[48][1] ),
    .ZN(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07213_ (.A1(\u2.mem[8][1] ),
    .A2(_02612_),
    .B1(_02614_),
    .B2(\u2.mem[4][1] ),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07214_ (.A1(\u2.mem[6][1] ),
    .A2(_02622_),
    .B1(_02624_),
    .B2(\u2.mem[47][1] ),
    .ZN(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07215_ (.A1(_02689_),
    .A2(_02690_),
    .A3(_02691_),
    .A4(_02692_),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07216_ (.A1(_02672_),
    .A2(_02679_),
    .A3(_02686_),
    .A4(_02693_),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07217_ (.A1(_01726_),
    .A2(_02361_),
    .B1(_02665_),
    .B2(_02694_),
    .ZN(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07218_ (.A1(\u2.mem[45][2] ),
    .A2(_02633_),
    .B1(_02634_),
    .B2(\u2.mem[34][2] ),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07219_ (.A1(\u2.mem[32][2] ),
    .A2(_02386_),
    .B1(_02396_),
    .B2(\u2.mem[2][2] ),
    .ZN(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07220_ (.A1(\u2.mem[40][2] ),
    .A2(_02406_),
    .B1(_02415_),
    .B2(\u2.mem[30][2] ),
    .ZN(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07221_ (.A1(\u2.mem[27][2] ),
    .A2(_02428_),
    .B1(_02436_),
    .B2(\u2.mem[35][2] ),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07222_ (.A1(_02695_),
    .A2(_02696_),
    .A3(_02697_),
    .A4(_02698_),
    .ZN(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07223_ (.A1(\u2.mem[15][2] ),
    .A2(_02457_),
    .B1(_02461_),
    .B2(\u2.mem[13][2] ),
    .ZN(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07224_ (.A1(\u2.mem[1][2] ),
    .A2(_02465_),
    .B1(_02471_),
    .B2(\u2.mem[7][2] ),
    .ZN(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07225_ (.A1(\u2.mem[16][2] ),
    .A2(_02475_),
    .B1(_02477_),
    .B2(\u2.mem[33][2] ),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07226_ (.A1(\u2.mem[3][2] ),
    .A2(_02480_),
    .B(_02359_),
    .ZN(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07227_ (.A1(_02700_),
    .A2(_02701_),
    .A3(_02702_),
    .A4(_02703_),
    .ZN(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07228_ (.A1(\u2.mem[50][2] ),
    .A2(_02645_),
    .B1(_02646_),
    .B2(\u2.mem[51][2] ),
    .ZN(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07229_ (.A1(\u2.mem[54][2] ),
    .A2(_02648_),
    .B1(_02649_),
    .B2(\u2.mem[55][2] ),
    .ZN(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07230_ (.A1(\u2.mem[53][2] ),
    .A2(_02486_),
    .B1(_02489_),
    .B2(\u2.mem[56][2] ),
    .ZN(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07231_ (.A1(\u2.mem[58][2] ),
    .A2(_02495_),
    .B1(_02500_),
    .B2(\u2.mem[36][2] ),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07232_ (.A1(_02705_),
    .A2(_02706_),
    .A3(_02707_),
    .A4(_02708_),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07233_ (.A1(\u2.mem[44][2] ),
    .A2(_02654_),
    .B1(_02655_),
    .B2(\u2.mem[42][2] ),
    .ZN(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07234_ (.A1(\u2.mem[14][2] ),
    .A2(_02657_),
    .B1(_02658_),
    .B2(\u2.mem[12][2] ),
    .ZN(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07235_ (.A1(\u2.mem[49][2] ),
    .A2(_02660_),
    .B1(_02661_),
    .B2(\u2.mem[46][2] ),
    .ZN(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07236_ (.A1(\u2.mem[43][2] ),
    .A2(_02515_),
    .B1(_02517_),
    .B2(\u2.mem[20][2] ),
    .ZN(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07237_ (.A1(_02710_),
    .A2(_02711_),
    .A3(_02712_),
    .A4(_02713_),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07238_ (.A1(_02699_),
    .A2(_02704_),
    .A3(_02709_),
    .A4(_02714_),
    .ZN(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07239_ (.A1(\u2.mem[61][2] ),
    .A2(_02666_),
    .B1(_02667_),
    .B2(\u2.mem[63][2] ),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07240_ (.A1(\u2.mem[60][2] ),
    .A2(_02546_),
    .B1(_02549_),
    .B2(\u2.mem[62][2] ),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07241_ (.A1(\u2.mem[37][2] ),
    .A2(_02540_),
    .B1(_02542_),
    .B2(\u2.mem[59][2] ),
    .ZN(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07242_ (.A1(\u2.mem[57][2] ),
    .A2(_02554_),
    .B1(_02556_),
    .B2(\u2.mem[41][2] ),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07243_ (.A1(_02716_),
    .A2(_02717_),
    .A3(_02718_),
    .A4(_02719_),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07244_ (.A1(\u2.mem[26][2] ),
    .A2(_02673_),
    .B1(_02674_),
    .B2(\u2.mem[10][2] ),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07245_ (.A1(\u2.mem[29][2] ),
    .A2(_02565_),
    .B1(_02570_),
    .B2(\u2.mem[11][2] ),
    .ZN(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07246_ (.A1(\u2.mem[9][2] ),
    .A2(_02580_),
    .B1(_02582_),
    .B2(\u2.mem[25][2] ),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07247_ (.A1(\u2.mem[28][2] ),
    .A2(_02585_),
    .B1(_02587_),
    .B2(\u2.mem[31][2] ),
    .ZN(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07248_ (.A1(_02721_),
    .A2(_02722_),
    .A3(_02723_),
    .A4(_02724_),
    .ZN(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07249_ (.A1(\u2.mem[23][2] ),
    .A2(_02680_),
    .B1(_02681_),
    .B2(\u2.mem[22][2] ),
    .ZN(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07250_ (.A1(\u2.mem[17][2] ),
    .A2(_02591_),
    .B1(_02593_),
    .B2(\u2.mem[24][2] ),
    .ZN(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07251_ (.A1(\u2.mem[52][2] ),
    .A2(_02601_),
    .B1(_02603_),
    .B2(\u2.mem[21][2] ),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07252_ (.A1(\u2.mem[18][2] ),
    .A2(_02606_),
    .B1(_02608_),
    .B2(\u2.mem[19][2] ),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07253_ (.A1(_02726_),
    .A2(_02727_),
    .A3(_02728_),
    .A4(_02729_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07254_ (.A1(\u2.mem[5][2] ),
    .A2(_02687_),
    .B1(_02688_),
    .B2(\u2.mem[38][2] ),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07255_ (.A1(\u2.mem[39][2] ),
    .A2(_02617_),
    .B1(_02619_),
    .B2(\u2.mem[48][2] ),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07256_ (.A1(\u2.mem[8][2] ),
    .A2(_02612_),
    .B1(_02614_),
    .B2(\u2.mem[4][2] ),
    .ZN(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07257_ (.A1(\u2.mem[6][2] ),
    .A2(_02622_),
    .B1(_02624_),
    .B2(\u2.mem[47][2] ),
    .ZN(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07258_ (.A1(_02731_),
    .A2(_02732_),
    .A3(_02733_),
    .A4(_02734_),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07259_ (.A1(_02720_),
    .A2(_02725_),
    .A3(_02730_),
    .A4(_02735_),
    .ZN(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07260_ (.A1(_01768_),
    .A2(_02361_),
    .B1(_02715_),
    .B2(_02736_),
    .ZN(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07261_ (.A1(\u2.mem[45][3] ),
    .A2(_02633_),
    .B1(_02634_),
    .B2(\u2.mem[34][3] ),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07262_ (.A1(\u2.mem[32][3] ),
    .A2(_02386_),
    .B1(_02396_),
    .B2(\u2.mem[2][3] ),
    .ZN(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07263_ (.A1(\u2.mem[40][3] ),
    .A2(_02406_),
    .B1(_02415_),
    .B2(\u2.mem[30][3] ),
    .ZN(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07264_ (.A1(\u2.mem[27][3] ),
    .A2(_02428_),
    .B1(_02436_),
    .B2(\u2.mem[35][3] ),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07265_ (.A1(_02737_),
    .A2(_02738_),
    .A3(_02739_),
    .A4(_02740_),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07266_ (.A1(\u2.mem[15][3] ),
    .A2(_02457_),
    .B1(_02461_),
    .B2(\u2.mem[13][3] ),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07267_ (.A1(\u2.mem[1][3] ),
    .A2(_02465_),
    .B1(_02471_),
    .B2(\u2.mem[7][3] ),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07268_ (.A1(\u2.mem[16][3] ),
    .A2(_02475_),
    .B1(_02477_),
    .B2(\u2.mem[33][3] ),
    .ZN(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07269_ (.I(_02358_),
    .Z(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07270_ (.A1(\u2.mem[3][3] ),
    .A2(_02480_),
    .B(_02745_),
    .ZN(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07271_ (.A1(_02742_),
    .A2(_02743_),
    .A3(_02744_),
    .A4(_02746_),
    .ZN(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07272_ (.A1(\u2.mem[50][3] ),
    .A2(_02645_),
    .B1(_02646_),
    .B2(\u2.mem[51][3] ),
    .ZN(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07273_ (.A1(\u2.mem[54][3] ),
    .A2(_02648_),
    .B1(_02649_),
    .B2(\u2.mem[55][3] ),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07274_ (.A1(\u2.mem[53][3] ),
    .A2(_02486_),
    .B1(_02489_),
    .B2(\u2.mem[56][3] ),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07275_ (.A1(\u2.mem[58][3] ),
    .A2(_02495_),
    .B1(_02500_),
    .B2(\u2.mem[36][3] ),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07276_ (.A1(_02748_),
    .A2(_02749_),
    .A3(_02750_),
    .A4(_02751_),
    .ZN(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07277_ (.A1(\u2.mem[44][3] ),
    .A2(_02654_),
    .B1(_02655_),
    .B2(\u2.mem[42][3] ),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07278_ (.A1(\u2.mem[14][3] ),
    .A2(_02657_),
    .B1(_02658_),
    .B2(\u2.mem[12][3] ),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07279_ (.A1(\u2.mem[49][3] ),
    .A2(_02660_),
    .B1(_02661_),
    .B2(\u2.mem[46][3] ),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07280_ (.A1(\u2.mem[43][3] ),
    .A2(_02515_),
    .B1(_02517_),
    .B2(\u2.mem[20][3] ),
    .ZN(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07281_ (.A1(_02753_),
    .A2(_02754_),
    .A3(_02755_),
    .A4(_02756_),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07282_ (.A1(_02741_),
    .A2(_02747_),
    .A3(_02752_),
    .A4(_02757_),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07283_ (.A1(\u2.mem[61][3] ),
    .A2(_02666_),
    .B1(_02667_),
    .B2(\u2.mem[63][3] ),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07284_ (.A1(\u2.mem[60][3] ),
    .A2(_02546_),
    .B1(_02549_),
    .B2(\u2.mem[62][3] ),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07285_ (.A1(\u2.mem[37][3] ),
    .A2(_02540_),
    .B1(_02542_),
    .B2(\u2.mem[59][3] ),
    .ZN(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07286_ (.A1(\u2.mem[57][3] ),
    .A2(_02554_),
    .B1(_02556_),
    .B2(\u2.mem[41][3] ),
    .ZN(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07287_ (.A1(_02759_),
    .A2(_02760_),
    .A3(_02761_),
    .A4(_02762_),
    .ZN(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07288_ (.A1(\u2.mem[26][3] ),
    .A2(_02673_),
    .B1(_02674_),
    .B2(\u2.mem[10][3] ),
    .ZN(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07289_ (.A1(\u2.mem[29][3] ),
    .A2(_02565_),
    .B1(_02570_),
    .B2(\u2.mem[11][3] ),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07290_ (.A1(\u2.mem[9][3] ),
    .A2(_02580_),
    .B1(_02582_),
    .B2(\u2.mem[25][3] ),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07291_ (.A1(\u2.mem[28][3] ),
    .A2(_02585_),
    .B1(_02587_),
    .B2(\u2.mem[31][3] ),
    .ZN(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07292_ (.A1(_02764_),
    .A2(_02765_),
    .A3(_02766_),
    .A4(_02767_),
    .ZN(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07293_ (.A1(\u2.mem[23][3] ),
    .A2(_02680_),
    .B1(_02681_),
    .B2(\u2.mem[22][3] ),
    .ZN(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07294_ (.A1(\u2.mem[17][3] ),
    .A2(_02591_),
    .B1(_02593_),
    .B2(\u2.mem[24][3] ),
    .ZN(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07295_ (.A1(\u2.mem[52][3] ),
    .A2(_02601_),
    .B1(_02603_),
    .B2(\u2.mem[21][3] ),
    .ZN(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07296_ (.A1(\u2.mem[18][3] ),
    .A2(_02606_),
    .B1(_02608_),
    .B2(\u2.mem[19][3] ),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07297_ (.A1(_02769_),
    .A2(_02770_),
    .A3(_02771_),
    .A4(_02772_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07298_ (.A1(\u2.mem[5][3] ),
    .A2(_02687_),
    .B1(_02688_),
    .B2(\u2.mem[38][3] ),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07299_ (.A1(\u2.mem[39][3] ),
    .A2(_02617_),
    .B1(_02619_),
    .B2(\u2.mem[48][3] ),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07300_ (.A1(\u2.mem[8][3] ),
    .A2(_02612_),
    .B1(_02614_),
    .B2(\u2.mem[4][3] ),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07301_ (.A1(\u2.mem[6][3] ),
    .A2(_02622_),
    .B1(_02624_),
    .B2(\u2.mem[47][3] ),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07302_ (.A1(_02774_),
    .A2(_02775_),
    .A3(_02776_),
    .A4(_02777_),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07303_ (.A1(_02763_),
    .A2(_02768_),
    .A3(_02773_),
    .A4(_02778_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07304_ (.A1(_01808_),
    .A2(_02361_),
    .B1(_02758_),
    .B2(_02779_),
    .ZN(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07305_ (.I(_02360_),
    .Z(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07306_ (.A1(\u2.mem[45][4] ),
    .A2(_02633_),
    .B1(_02634_),
    .B2(\u2.mem[34][4] ),
    .ZN(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07307_ (.I(_02385_),
    .Z(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07308_ (.I(_02395_),
    .Z(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07309_ (.A1(\u2.mem[32][4] ),
    .A2(_02782_),
    .B1(_02783_),
    .B2(\u2.mem[2][4] ),
    .ZN(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07310_ (.I(_02405_),
    .Z(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07311_ (.I(_02414_),
    .Z(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07312_ (.A1(\u2.mem[40][4] ),
    .A2(_02785_),
    .B1(_02786_),
    .B2(\u2.mem[30][4] ),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07313_ (.I(_02427_),
    .Z(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07314_ (.I(_02435_),
    .Z(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07315_ (.A1(\u2.mem[27][4] ),
    .A2(_02788_),
    .B1(_02789_),
    .B2(\u2.mem[35][4] ),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07316_ (.A1(_02781_),
    .A2(_02784_),
    .A3(_02787_),
    .A4(_02790_),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07317_ (.I(_02456_),
    .Z(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07318_ (.I(_02460_),
    .Z(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07319_ (.A1(\u2.mem[15][4] ),
    .A2(_02792_),
    .B1(_02793_),
    .B2(\u2.mem[13][4] ),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07320_ (.I(_02464_),
    .Z(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07321_ (.I(_02470_),
    .Z(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07322_ (.A1(\u2.mem[1][4] ),
    .A2(_02795_),
    .B1(_02796_),
    .B2(\u2.mem[7][4] ),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07323_ (.I(_02474_),
    .Z(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07324_ (.I(_02476_),
    .Z(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07325_ (.A1(\u2.mem[16][4] ),
    .A2(_02798_),
    .B1(_02799_),
    .B2(\u2.mem[33][4] ),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07326_ (.I(_02479_),
    .Z(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07327_ (.A1(\u2.mem[3][4] ),
    .A2(_02801_),
    .B(_02745_),
    .ZN(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07328_ (.A1(_02794_),
    .A2(_02797_),
    .A3(_02800_),
    .A4(_02802_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07329_ (.A1(\u2.mem[50][4] ),
    .A2(_02645_),
    .B1(_02646_),
    .B2(\u2.mem[51][4] ),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07330_ (.A1(\u2.mem[54][4] ),
    .A2(_02648_),
    .B1(_02649_),
    .B2(\u2.mem[55][4] ),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07331_ (.I(_02485_),
    .Z(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07332_ (.I(_02488_),
    .Z(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07333_ (.A1(\u2.mem[53][4] ),
    .A2(_02806_),
    .B1(_02807_),
    .B2(\u2.mem[56][4] ),
    .ZN(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07334_ (.I(_02494_),
    .Z(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07335_ (.I(_02499_),
    .Z(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07336_ (.A1(\u2.mem[58][4] ),
    .A2(_02809_),
    .B1(_02810_),
    .B2(\u2.mem[36][4] ),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07337_ (.A1(_02804_),
    .A2(_02805_),
    .A3(_02808_),
    .A4(_02811_),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07338_ (.A1(\u2.mem[44][4] ),
    .A2(_02654_),
    .B1(_02655_),
    .B2(\u2.mem[42][4] ),
    .ZN(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07339_ (.A1(\u2.mem[14][4] ),
    .A2(_02657_),
    .B1(_02658_),
    .B2(\u2.mem[12][4] ),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07340_ (.A1(\u2.mem[49][4] ),
    .A2(_02660_),
    .B1(_02661_),
    .B2(\u2.mem[46][4] ),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07341_ (.I(_02514_),
    .Z(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07342_ (.I(_02516_),
    .Z(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07343_ (.A1(\u2.mem[43][4] ),
    .A2(_02816_),
    .B1(_02817_),
    .B2(\u2.mem[20][4] ),
    .ZN(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07344_ (.A1(_02813_),
    .A2(_02814_),
    .A3(_02815_),
    .A4(_02818_),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07345_ (.A1(_02791_),
    .A2(_02803_),
    .A3(_02812_),
    .A4(_02819_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07346_ (.A1(\u2.mem[61][4] ),
    .A2(_02666_),
    .B1(_02667_),
    .B2(\u2.mem[63][4] ),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07347_ (.I(_02545_),
    .Z(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07348_ (.I(_02548_),
    .Z(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07349_ (.A1(\u2.mem[60][4] ),
    .A2(_02822_),
    .B1(_02823_),
    .B2(\u2.mem[62][4] ),
    .ZN(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07350_ (.I(_02539_),
    .Z(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07351_ (.I(_02541_),
    .Z(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07352_ (.A1(\u2.mem[37][4] ),
    .A2(_02825_),
    .B1(_02826_),
    .B2(\u2.mem[59][4] ),
    .ZN(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07353_ (.I(_02553_),
    .Z(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07354_ (.I(_02555_),
    .Z(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07355_ (.A1(\u2.mem[57][4] ),
    .A2(_02828_),
    .B1(_02829_),
    .B2(\u2.mem[41][4] ),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07356_ (.A1(_02821_),
    .A2(_02824_),
    .A3(_02827_),
    .A4(_02830_),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07357_ (.A1(\u2.mem[26][4] ),
    .A2(_02673_),
    .B1(_02674_),
    .B2(\u2.mem[10][4] ),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07358_ (.I(_02564_),
    .Z(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07359_ (.I(_02569_),
    .Z(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07360_ (.A1(\u2.mem[29][4] ),
    .A2(_02833_),
    .B1(_02834_),
    .B2(\u2.mem[11][4] ),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07361_ (.I(_02579_),
    .Z(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07362_ (.I(_02581_),
    .Z(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07363_ (.A1(\u2.mem[9][4] ),
    .A2(_02836_),
    .B1(_02837_),
    .B2(\u2.mem[25][4] ),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07364_ (.I(_02584_),
    .Z(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07365_ (.I(_02586_),
    .Z(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07366_ (.A1(\u2.mem[28][4] ),
    .A2(_02839_),
    .B1(_02840_),
    .B2(\u2.mem[31][4] ),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07367_ (.A1(_02832_),
    .A2(_02835_),
    .A3(_02838_),
    .A4(_02841_),
    .ZN(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07368_ (.A1(\u2.mem[23][4] ),
    .A2(_02680_),
    .B1(_02681_),
    .B2(\u2.mem[22][4] ),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07369_ (.I(_02590_),
    .Z(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07370_ (.I(_02592_),
    .Z(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07371_ (.A1(\u2.mem[17][4] ),
    .A2(_02844_),
    .B1(_02845_),
    .B2(\u2.mem[24][4] ),
    .ZN(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07372_ (.I(_02600_),
    .Z(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07373_ (.I(_02602_),
    .Z(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07374_ (.A1(\u2.mem[52][4] ),
    .A2(_02847_),
    .B1(_02848_),
    .B2(\u2.mem[21][4] ),
    .ZN(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07375_ (.I(_02605_),
    .Z(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07376_ (.I(_02607_),
    .Z(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07377_ (.A1(\u2.mem[18][4] ),
    .A2(_02850_),
    .B1(_02851_),
    .B2(\u2.mem[19][4] ),
    .ZN(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07378_ (.A1(_02843_),
    .A2(_02846_),
    .A3(_02849_),
    .A4(_02852_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07379_ (.A1(\u2.mem[5][4] ),
    .A2(_02687_),
    .B1(_02688_),
    .B2(\u2.mem[38][4] ),
    .ZN(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07380_ (.I(_02616_),
    .Z(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07381_ (.I(_02618_),
    .Z(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07382_ (.A1(\u2.mem[39][4] ),
    .A2(_02855_),
    .B1(_02856_),
    .B2(\u2.mem[48][4] ),
    .ZN(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07383_ (.I(_02611_),
    .Z(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07384_ (.I(_02613_),
    .Z(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07385_ (.A1(\u2.mem[8][4] ),
    .A2(_02858_),
    .B1(_02859_),
    .B2(\u2.mem[4][4] ),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07386_ (.I(_02621_),
    .Z(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07387_ (.I(_02623_),
    .Z(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07388_ (.A1(\u2.mem[6][4] ),
    .A2(_02861_),
    .B1(_02862_),
    .B2(\u2.mem[47][4] ),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07389_ (.A1(_02854_),
    .A2(_02857_),
    .A3(_02860_),
    .A4(_02863_),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07390_ (.A1(_02831_),
    .A2(_02842_),
    .A3(_02853_),
    .A4(_02864_),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07391_ (.A1(_01843_),
    .A2(_02780_),
    .B1(_02820_),
    .B2(_02865_),
    .ZN(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07392_ (.I(_02443_),
    .Z(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07393_ (.I(_02447_),
    .Z(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07394_ (.A1(\u2.mem[45][5] ),
    .A2(_02866_),
    .B1(_02867_),
    .B2(\u2.mem[34][5] ),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07395_ (.A1(\u2.mem[32][5] ),
    .A2(_02782_),
    .B1(_02783_),
    .B2(\u2.mem[2][5] ),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07396_ (.A1(\u2.mem[40][5] ),
    .A2(_02785_),
    .B1(_02786_),
    .B2(\u2.mem[30][5] ),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07397_ (.A1(\u2.mem[27][5] ),
    .A2(_02788_),
    .B1(_02789_),
    .B2(\u2.mem[35][5] ),
    .ZN(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07398_ (.A1(_02868_),
    .A2(_02869_),
    .A3(_02870_),
    .A4(_02871_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07399_ (.A1(\u2.mem[15][5] ),
    .A2(_02792_),
    .B1(_02793_),
    .B2(\u2.mem[13][5] ),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07400_ (.A1(\u2.mem[1][5] ),
    .A2(_02795_),
    .B1(_02796_),
    .B2(\u2.mem[7][5] ),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07401_ (.A1(\u2.mem[16][5] ),
    .A2(_02798_),
    .B1(_02799_),
    .B2(\u2.mem[33][5] ),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07402_ (.A1(\u2.mem[3][5] ),
    .A2(_02801_),
    .B(_02745_),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07403_ (.A1(_02873_),
    .A2(_02874_),
    .A3(_02875_),
    .A4(_02876_),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07404_ (.I(_02502_),
    .Z(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07405_ (.I(_02504_),
    .Z(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07406_ (.A1(\u2.mem[50][5] ),
    .A2(_02878_),
    .B1(_02879_),
    .B2(\u2.mem[51][5] ),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07407_ (.I(_02508_),
    .Z(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07408_ (.I(_02510_),
    .Z(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07409_ (.A1(\u2.mem[54][5] ),
    .A2(_02881_),
    .B1(_02882_),
    .B2(\u2.mem[55][5] ),
    .ZN(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07410_ (.A1(\u2.mem[53][5] ),
    .A2(_02806_),
    .B1(_02807_),
    .B2(\u2.mem[56][5] ),
    .ZN(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07411_ (.A1(\u2.mem[58][5] ),
    .A2(_02809_),
    .B1(_02810_),
    .B2(\u2.mem[36][5] ),
    .ZN(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07412_ (.A1(_02880_),
    .A2(_02883_),
    .A3(_02884_),
    .A4(_02885_),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07413_ (.I(_02520_),
    .Z(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07414_ (.I(_02522_),
    .Z(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07415_ (.A1(\u2.mem[44][5] ),
    .A2(_02887_),
    .B1(_02888_),
    .B2(\u2.mem[42][5] ),
    .ZN(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07416_ (.I(_02525_),
    .Z(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07417_ (.I(_02527_),
    .Z(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07418_ (.A1(\u2.mem[14][5] ),
    .A2(_02890_),
    .B1(_02891_),
    .B2(\u2.mem[12][5] ),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07419_ (.I(_02530_),
    .Z(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07420_ (.I(_02532_),
    .Z(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07421_ (.A1(\u2.mem[49][5] ),
    .A2(_02893_),
    .B1(_02894_),
    .B2(\u2.mem[46][5] ),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07422_ (.A1(\u2.mem[43][5] ),
    .A2(_02816_),
    .B1(_02817_),
    .B2(\u2.mem[20][5] ),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07423_ (.A1(_02889_),
    .A2(_02892_),
    .A3(_02895_),
    .A4(_02896_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07424_ (.A1(_02872_),
    .A2(_02877_),
    .A3(_02886_),
    .A4(_02897_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07425_ (.I(_02558_),
    .Z(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07426_ (.I(_02560_),
    .Z(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07427_ (.A1(\u2.mem[61][5] ),
    .A2(_02899_),
    .B1(_02900_),
    .B2(\u2.mem[63][5] ),
    .ZN(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07428_ (.A1(\u2.mem[60][5] ),
    .A2(_02822_),
    .B1(_02823_),
    .B2(\u2.mem[62][5] ),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07429_ (.A1(\u2.mem[37][5] ),
    .A2(_02825_),
    .B1(_02826_),
    .B2(\u2.mem[59][5] ),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07430_ (.A1(\u2.mem[57][5] ),
    .A2(_02828_),
    .B1(_02829_),
    .B2(\u2.mem[41][5] ),
    .ZN(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07431_ (.A1(_02901_),
    .A2(_02902_),
    .A3(_02903_),
    .A4(_02904_),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07432_ (.I(_02572_),
    .Z(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07433_ (.I(_02574_),
    .Z(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07434_ (.A1(\u2.mem[26][5] ),
    .A2(_02906_),
    .B1(_02907_),
    .B2(\u2.mem[10][5] ),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07435_ (.A1(\u2.mem[29][5] ),
    .A2(_02833_),
    .B1(_02834_),
    .B2(\u2.mem[11][5] ),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07436_ (.A1(\u2.mem[9][5] ),
    .A2(_02836_),
    .B1(_02837_),
    .B2(\u2.mem[25][5] ),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07437_ (.A1(\u2.mem[28][5] ),
    .A2(_02839_),
    .B1(_02840_),
    .B2(\u2.mem[31][5] ),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07438_ (.A1(_02908_),
    .A2(_02909_),
    .A3(_02910_),
    .A4(_02911_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07439_ (.I(_02595_),
    .Z(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07440_ (.I(_02597_),
    .Z(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07441_ (.A1(\u2.mem[23][5] ),
    .A2(_02913_),
    .B1(_02914_),
    .B2(\u2.mem[22][5] ),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07442_ (.A1(\u2.mem[17][5] ),
    .A2(_02844_),
    .B1(_02845_),
    .B2(\u2.mem[24][5] ),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07443_ (.A1(\u2.mem[52][5] ),
    .A2(_02847_),
    .B1(_02848_),
    .B2(\u2.mem[21][5] ),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07444_ (.A1(\u2.mem[18][5] ),
    .A2(_02850_),
    .B1(_02851_),
    .B2(\u2.mem[19][5] ),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07445_ (.A1(_02915_),
    .A2(_02916_),
    .A3(_02917_),
    .A4(_02918_),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07446_ (.I(_02626_),
    .Z(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07447_ (.I(_02628_),
    .Z(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07448_ (.A1(\u2.mem[5][5] ),
    .A2(_02920_),
    .B1(_02921_),
    .B2(\u2.mem[38][5] ),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07449_ (.A1(\u2.mem[39][5] ),
    .A2(_02855_),
    .B1(_02856_),
    .B2(\u2.mem[48][5] ),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07450_ (.A1(\u2.mem[8][5] ),
    .A2(_02858_),
    .B1(_02859_),
    .B2(\u2.mem[4][5] ),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07451_ (.A1(\u2.mem[6][5] ),
    .A2(_02861_),
    .B1(_02862_),
    .B2(\u2.mem[47][5] ),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07452_ (.A1(_02922_),
    .A2(_02923_),
    .A3(_02924_),
    .A4(_02925_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07453_ (.A1(_02905_),
    .A2(_02912_),
    .A3(_02919_),
    .A4(_02926_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07454_ (.A1(_01877_),
    .A2(_02780_),
    .B1(_02898_),
    .B2(_02927_),
    .ZN(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07455_ (.A1(\u2.mem[45][6] ),
    .A2(_02866_),
    .B1(_02867_),
    .B2(\u2.mem[34][6] ),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07456_ (.A1(\u2.mem[32][6] ),
    .A2(_02782_),
    .B1(_02783_),
    .B2(\u2.mem[2][6] ),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07457_ (.A1(\u2.mem[40][6] ),
    .A2(_02785_),
    .B1(_02786_),
    .B2(\u2.mem[30][6] ),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07458_ (.A1(\u2.mem[27][6] ),
    .A2(_02788_),
    .B1(_02789_),
    .B2(\u2.mem[35][6] ),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07459_ (.A1(_02928_),
    .A2(_02929_),
    .A3(_02930_),
    .A4(_02931_),
    .ZN(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07460_ (.A1(\u2.mem[15][6] ),
    .A2(_02792_),
    .B1(_02793_),
    .B2(\u2.mem[13][6] ),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07461_ (.A1(\u2.mem[1][6] ),
    .A2(_02795_),
    .B1(_02796_),
    .B2(\u2.mem[7][6] ),
    .ZN(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07462_ (.A1(\u2.mem[16][6] ),
    .A2(_02798_),
    .B1(_02799_),
    .B2(\u2.mem[33][6] ),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07463_ (.A1(\u2.mem[3][6] ),
    .A2(_02801_),
    .B(_02745_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07464_ (.A1(_02933_),
    .A2(_02934_),
    .A3(_02935_),
    .A4(_02936_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07465_ (.A1(\u2.mem[50][6] ),
    .A2(_02878_),
    .B1(_02879_),
    .B2(\u2.mem[51][6] ),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07466_ (.A1(\u2.mem[54][6] ),
    .A2(_02881_),
    .B1(_02882_),
    .B2(\u2.mem[55][6] ),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07467_ (.A1(\u2.mem[53][6] ),
    .A2(_02806_),
    .B1(_02807_),
    .B2(\u2.mem[56][6] ),
    .ZN(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07468_ (.A1(\u2.mem[58][6] ),
    .A2(_02809_),
    .B1(_02810_),
    .B2(\u2.mem[36][6] ),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07469_ (.A1(_02938_),
    .A2(_02939_),
    .A3(_02940_),
    .A4(_02941_),
    .ZN(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07470_ (.A1(\u2.mem[44][6] ),
    .A2(_02887_),
    .B1(_02888_),
    .B2(\u2.mem[42][6] ),
    .ZN(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07471_ (.A1(\u2.mem[14][6] ),
    .A2(_02890_),
    .B1(_02891_),
    .B2(\u2.mem[12][6] ),
    .ZN(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07472_ (.A1(\u2.mem[49][6] ),
    .A2(_02893_),
    .B1(_02894_),
    .B2(\u2.mem[46][6] ),
    .ZN(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07473_ (.A1(\u2.mem[43][6] ),
    .A2(_02816_),
    .B1(_02817_),
    .B2(\u2.mem[20][6] ),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07474_ (.A1(_02943_),
    .A2(_02944_),
    .A3(_02945_),
    .A4(_02946_),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07475_ (.A1(_02932_),
    .A2(_02937_),
    .A3(_02942_),
    .A4(_02947_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07476_ (.A1(\u2.mem[61][6] ),
    .A2(_02899_),
    .B1(_02900_),
    .B2(\u2.mem[63][6] ),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07477_ (.A1(\u2.mem[60][6] ),
    .A2(_02822_),
    .B1(_02823_),
    .B2(\u2.mem[62][6] ),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07478_ (.A1(\u2.mem[37][6] ),
    .A2(_02825_),
    .B1(_02826_),
    .B2(\u2.mem[59][6] ),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07479_ (.A1(\u2.mem[57][6] ),
    .A2(_02828_),
    .B1(_02829_),
    .B2(\u2.mem[41][6] ),
    .ZN(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07480_ (.A1(_02949_),
    .A2(_02950_),
    .A3(_02951_),
    .A4(_02952_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07481_ (.A1(\u2.mem[26][6] ),
    .A2(_02906_),
    .B1(_02907_),
    .B2(\u2.mem[10][6] ),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07482_ (.A1(\u2.mem[29][6] ),
    .A2(_02833_),
    .B1(_02834_),
    .B2(\u2.mem[11][6] ),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07483_ (.A1(\u2.mem[9][6] ),
    .A2(_02836_),
    .B1(_02837_),
    .B2(\u2.mem[25][6] ),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07484_ (.A1(\u2.mem[28][6] ),
    .A2(_02839_),
    .B1(_02840_),
    .B2(\u2.mem[31][6] ),
    .ZN(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07485_ (.A1(_02954_),
    .A2(_02955_),
    .A3(_02956_),
    .A4(_02957_),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07486_ (.A1(\u2.mem[23][6] ),
    .A2(_02913_),
    .B1(_02914_),
    .B2(\u2.mem[22][6] ),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07487_ (.A1(\u2.mem[17][6] ),
    .A2(_02844_),
    .B1(_02845_),
    .B2(\u2.mem[24][6] ),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07488_ (.A1(\u2.mem[52][6] ),
    .A2(_02847_),
    .B1(_02848_),
    .B2(\u2.mem[21][6] ),
    .ZN(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07489_ (.A1(\u2.mem[18][6] ),
    .A2(_02850_),
    .B1(_02851_),
    .B2(\u2.mem[19][6] ),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07490_ (.A1(_02959_),
    .A2(_02960_),
    .A3(_02961_),
    .A4(_02962_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07491_ (.A1(\u2.mem[5][6] ),
    .A2(_02920_),
    .B1(_02921_),
    .B2(\u2.mem[38][6] ),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07492_ (.A1(\u2.mem[39][6] ),
    .A2(_02855_),
    .B1(_02856_),
    .B2(\u2.mem[48][6] ),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07493_ (.A1(\u2.mem[8][6] ),
    .A2(_02858_),
    .B1(_02859_),
    .B2(\u2.mem[4][6] ),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07494_ (.A1(\u2.mem[6][6] ),
    .A2(_02861_),
    .B1(_02862_),
    .B2(\u2.mem[47][6] ),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07495_ (.A1(_02964_),
    .A2(_02965_),
    .A3(_02966_),
    .A4(_02967_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07496_ (.A1(_02953_),
    .A2(_02958_),
    .A3(_02963_),
    .A4(_02968_),
    .ZN(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07497_ (.A1(_01945_),
    .A2(_02780_),
    .B1(_02948_),
    .B2(_02969_),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07498_ (.A1(\u2.mem[45][7] ),
    .A2(_02866_),
    .B1(_02867_),
    .B2(\u2.mem[34][7] ),
    .ZN(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07499_ (.A1(\u2.mem[32][7] ),
    .A2(_02782_),
    .B1(_02783_),
    .B2(\u2.mem[2][7] ),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07500_ (.A1(\u2.mem[40][7] ),
    .A2(_02785_),
    .B1(_02786_),
    .B2(\u2.mem[30][7] ),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07501_ (.A1(\u2.mem[27][7] ),
    .A2(_02788_),
    .B1(_02789_),
    .B2(\u2.mem[35][7] ),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07502_ (.A1(_02970_),
    .A2(_02971_),
    .A3(_02972_),
    .A4(_02973_),
    .ZN(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07503_ (.A1(\u2.mem[15][7] ),
    .A2(_02792_),
    .B1(_02793_),
    .B2(\u2.mem[13][7] ),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07504_ (.A1(\u2.mem[1][7] ),
    .A2(_02795_),
    .B1(_02796_),
    .B2(\u2.mem[7][7] ),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07505_ (.A1(\u2.mem[16][7] ),
    .A2(_02798_),
    .B1(_02799_),
    .B2(\u2.mem[33][7] ),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07506_ (.I(_02358_),
    .Z(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07507_ (.A1(\u2.mem[3][7] ),
    .A2(_02801_),
    .B(_02978_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07508_ (.A1(_02975_),
    .A2(_02976_),
    .A3(_02977_),
    .A4(_02979_),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07509_ (.A1(\u2.mem[50][7] ),
    .A2(_02878_),
    .B1(_02879_),
    .B2(\u2.mem[51][7] ),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07510_ (.A1(\u2.mem[54][7] ),
    .A2(_02881_),
    .B1(_02882_),
    .B2(\u2.mem[55][7] ),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07511_ (.A1(\u2.mem[53][7] ),
    .A2(_02806_),
    .B1(_02807_),
    .B2(\u2.mem[56][7] ),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07512_ (.A1(\u2.mem[58][7] ),
    .A2(_02809_),
    .B1(_02810_),
    .B2(\u2.mem[36][7] ),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07513_ (.A1(_02981_),
    .A2(_02982_),
    .A3(_02983_),
    .A4(_02984_),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07514_ (.A1(\u2.mem[44][7] ),
    .A2(_02887_),
    .B1(_02888_),
    .B2(\u2.mem[42][7] ),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07515_ (.A1(\u2.mem[14][7] ),
    .A2(_02890_),
    .B1(_02891_),
    .B2(\u2.mem[12][7] ),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07516_ (.A1(\u2.mem[49][7] ),
    .A2(_02893_),
    .B1(_02894_),
    .B2(\u2.mem[46][7] ),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07517_ (.A1(\u2.mem[43][7] ),
    .A2(_02816_),
    .B1(_02817_),
    .B2(\u2.mem[20][7] ),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07518_ (.A1(_02986_),
    .A2(_02987_),
    .A3(_02988_),
    .A4(_02989_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07519_ (.A1(_02974_),
    .A2(_02980_),
    .A3(_02985_),
    .A4(_02990_),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07520_ (.A1(\u2.mem[61][7] ),
    .A2(_02899_),
    .B1(_02900_),
    .B2(\u2.mem[63][7] ),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07521_ (.A1(\u2.mem[60][7] ),
    .A2(_02822_),
    .B1(_02823_),
    .B2(\u2.mem[62][7] ),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07522_ (.A1(\u2.mem[37][7] ),
    .A2(_02825_),
    .B1(_02826_),
    .B2(\u2.mem[59][7] ),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07523_ (.A1(\u2.mem[57][7] ),
    .A2(_02828_),
    .B1(_02829_),
    .B2(\u2.mem[41][7] ),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07524_ (.A1(_02992_),
    .A2(_02993_),
    .A3(_02994_),
    .A4(_02995_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07525_ (.A1(\u2.mem[26][7] ),
    .A2(_02906_),
    .B1(_02907_),
    .B2(\u2.mem[10][7] ),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07526_ (.A1(\u2.mem[29][7] ),
    .A2(_02833_),
    .B1(_02834_),
    .B2(\u2.mem[11][7] ),
    .ZN(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07527_ (.A1(\u2.mem[9][7] ),
    .A2(_02836_),
    .B1(_02837_),
    .B2(\u2.mem[25][7] ),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07528_ (.A1(\u2.mem[28][7] ),
    .A2(_02839_),
    .B1(_02840_),
    .B2(\u2.mem[31][7] ),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07529_ (.A1(_02997_),
    .A2(_02998_),
    .A3(_02999_),
    .A4(_03000_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07530_ (.A1(\u2.mem[23][7] ),
    .A2(_02913_),
    .B1(_02914_),
    .B2(\u2.mem[22][7] ),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07531_ (.A1(\u2.mem[17][7] ),
    .A2(_02844_),
    .B1(_02845_),
    .B2(\u2.mem[24][7] ),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07532_ (.A1(\u2.mem[52][7] ),
    .A2(_02847_),
    .B1(_02848_),
    .B2(\u2.mem[21][7] ),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07533_ (.A1(\u2.mem[18][7] ),
    .A2(_02850_),
    .B1(_02851_),
    .B2(\u2.mem[19][7] ),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07534_ (.A1(_03002_),
    .A2(_03003_),
    .A3(_03004_),
    .A4(_03005_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07535_ (.A1(\u2.mem[5][7] ),
    .A2(_02920_),
    .B1(_02921_),
    .B2(\u2.mem[38][7] ),
    .ZN(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07536_ (.A1(\u2.mem[39][7] ),
    .A2(_02855_),
    .B1(_02856_),
    .B2(\u2.mem[48][7] ),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07537_ (.A1(\u2.mem[8][7] ),
    .A2(_02858_),
    .B1(_02859_),
    .B2(\u2.mem[4][7] ),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07538_ (.A1(\u2.mem[6][7] ),
    .A2(_02861_),
    .B1(_02862_),
    .B2(\u2.mem[47][7] ),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07539_ (.A1(_03007_),
    .A2(_03008_),
    .A3(_03009_),
    .A4(_03010_),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07540_ (.A1(_02996_),
    .A2(_03001_),
    .A3(_03006_),
    .A4(_03011_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07541_ (.A1(_01951_),
    .A2(_02780_),
    .B1(_02991_),
    .B2(_03012_),
    .ZN(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07542_ (.I(_02360_),
    .Z(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07543_ (.A1(\u2.mem[45][8] ),
    .A2(_02866_),
    .B1(_02867_),
    .B2(\u2.mem[34][8] ),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07544_ (.I(_02385_),
    .Z(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07545_ (.I(_02395_),
    .Z(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07546_ (.A1(\u2.mem[32][8] ),
    .A2(_03015_),
    .B1(_03016_),
    .B2(\u2.mem[2][8] ),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07547_ (.I(_02405_),
    .Z(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07548_ (.I(_02414_),
    .Z(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07549_ (.A1(\u2.mem[40][8] ),
    .A2(_03018_),
    .B1(_03019_),
    .B2(\u2.mem[30][8] ),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07550_ (.I(_02427_),
    .Z(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07551_ (.I(_02435_),
    .Z(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07552_ (.A1(\u2.mem[27][8] ),
    .A2(_03021_),
    .B1(_03022_),
    .B2(\u2.mem[35][8] ),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07553_ (.A1(_03014_),
    .A2(_03017_),
    .A3(_03020_),
    .A4(_03023_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07554_ (.I(_02456_),
    .Z(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07555_ (.I(_02460_),
    .Z(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07556_ (.A1(\u2.mem[15][8] ),
    .A2(_03025_),
    .B1(_03026_),
    .B2(\u2.mem[13][8] ),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07557_ (.I(_02464_),
    .Z(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07558_ (.I(_02470_),
    .Z(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07559_ (.A1(\u2.mem[1][8] ),
    .A2(_03028_),
    .B1(_03029_),
    .B2(\u2.mem[7][8] ),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07560_ (.I(_02474_),
    .Z(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07561_ (.I(_02476_),
    .Z(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07562_ (.A1(\u2.mem[16][8] ),
    .A2(_03031_),
    .B1(_03032_),
    .B2(\u2.mem[33][8] ),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07563_ (.I(_02479_),
    .Z(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07564_ (.A1(\u2.mem[3][8] ),
    .A2(_03034_),
    .B(_02978_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07565_ (.A1(_03027_),
    .A2(_03030_),
    .A3(_03033_),
    .A4(_03035_),
    .ZN(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07566_ (.A1(\u2.mem[50][8] ),
    .A2(_02878_),
    .B1(_02879_),
    .B2(\u2.mem[51][8] ),
    .ZN(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07567_ (.A1(\u2.mem[54][8] ),
    .A2(_02881_),
    .B1(_02882_),
    .B2(\u2.mem[55][8] ),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07568_ (.I(_02485_),
    .Z(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07569_ (.I(_02488_),
    .Z(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07570_ (.A1(\u2.mem[53][8] ),
    .A2(_03039_),
    .B1(_03040_),
    .B2(\u2.mem[56][8] ),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07571_ (.I(_02494_),
    .Z(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07572_ (.I(_02499_),
    .Z(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07573_ (.A1(\u2.mem[58][8] ),
    .A2(_03042_),
    .B1(_03043_),
    .B2(\u2.mem[36][8] ),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07574_ (.A1(_03037_),
    .A2(_03038_),
    .A3(_03041_),
    .A4(_03044_),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07575_ (.A1(\u2.mem[44][8] ),
    .A2(_02887_),
    .B1(_02888_),
    .B2(\u2.mem[42][8] ),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07576_ (.A1(\u2.mem[14][8] ),
    .A2(_02890_),
    .B1(_02891_),
    .B2(\u2.mem[12][8] ),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07577_ (.A1(\u2.mem[49][8] ),
    .A2(_02893_),
    .B1(_02894_),
    .B2(\u2.mem[46][8] ),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07578_ (.I(_02514_),
    .Z(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07579_ (.I(_02516_),
    .Z(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07580_ (.A1(\u2.mem[43][8] ),
    .A2(_03049_),
    .B1(_03050_),
    .B2(\u2.mem[20][8] ),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07581_ (.A1(_03046_),
    .A2(_03047_),
    .A3(_03048_),
    .A4(_03051_),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07582_ (.A1(_03024_),
    .A2(_03036_),
    .A3(_03045_),
    .A4(_03052_),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07583_ (.A1(\u2.mem[61][8] ),
    .A2(_02899_),
    .B1(_02900_),
    .B2(\u2.mem[63][8] ),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07584_ (.I(_02545_),
    .Z(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07585_ (.I(_02548_),
    .Z(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07586_ (.A1(\u2.mem[60][8] ),
    .A2(_03055_),
    .B1(_03056_),
    .B2(\u2.mem[62][8] ),
    .ZN(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07587_ (.I(_02539_),
    .Z(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07588_ (.I(_02541_),
    .Z(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07589_ (.A1(\u2.mem[37][8] ),
    .A2(_03058_),
    .B1(_03059_),
    .B2(\u2.mem[59][8] ),
    .ZN(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07590_ (.I(_02553_),
    .Z(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07591_ (.I(_02555_),
    .Z(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07592_ (.A1(\u2.mem[57][8] ),
    .A2(_03061_),
    .B1(_03062_),
    .B2(\u2.mem[41][8] ),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07593_ (.A1(_03054_),
    .A2(_03057_),
    .A3(_03060_),
    .A4(_03063_),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07594_ (.A1(\u2.mem[26][8] ),
    .A2(_02906_),
    .B1(_02907_),
    .B2(\u2.mem[10][8] ),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07595_ (.I(_02564_),
    .Z(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07596_ (.I(_02569_),
    .Z(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07597_ (.A1(\u2.mem[29][8] ),
    .A2(_03066_),
    .B1(_03067_),
    .B2(\u2.mem[11][8] ),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07598_ (.I(_02579_),
    .Z(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07599_ (.I(_02581_),
    .Z(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07600_ (.A1(\u2.mem[9][8] ),
    .A2(_03069_),
    .B1(_03070_),
    .B2(\u2.mem[25][8] ),
    .ZN(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07601_ (.I(_02584_),
    .Z(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07602_ (.I(_02586_),
    .Z(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07603_ (.A1(\u2.mem[28][8] ),
    .A2(_03072_),
    .B1(_03073_),
    .B2(\u2.mem[31][8] ),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07604_ (.A1(_03065_),
    .A2(_03068_),
    .A3(_03071_),
    .A4(_03074_),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07605_ (.A1(\u2.mem[23][8] ),
    .A2(_02913_),
    .B1(_02914_),
    .B2(\u2.mem[22][8] ),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07606_ (.I(_02590_),
    .Z(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07607_ (.I(_02592_),
    .Z(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07608_ (.A1(\u2.mem[17][8] ),
    .A2(_03077_),
    .B1(_03078_),
    .B2(\u2.mem[24][8] ),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07609_ (.I(_02600_),
    .Z(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07610_ (.I(_02602_),
    .Z(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07611_ (.A1(\u2.mem[52][8] ),
    .A2(_03080_),
    .B1(_03081_),
    .B2(\u2.mem[21][8] ),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07612_ (.I(_02605_),
    .Z(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07613_ (.I(_02607_),
    .Z(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07614_ (.A1(\u2.mem[18][8] ),
    .A2(_03083_),
    .B1(_03084_),
    .B2(\u2.mem[19][8] ),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07615_ (.A1(_03076_),
    .A2(_03079_),
    .A3(_03082_),
    .A4(_03085_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07616_ (.A1(\u2.mem[5][8] ),
    .A2(_02920_),
    .B1(_02921_),
    .B2(\u2.mem[38][8] ),
    .ZN(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07617_ (.I(_02616_),
    .Z(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07618_ (.I(_02618_),
    .Z(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07619_ (.A1(\u2.mem[39][8] ),
    .A2(_03088_),
    .B1(_03089_),
    .B2(\u2.mem[48][8] ),
    .ZN(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07620_ (.I(_02611_),
    .Z(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07621_ (.I(_02613_),
    .Z(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07622_ (.A1(\u2.mem[8][8] ),
    .A2(_03091_),
    .B1(_03092_),
    .B2(\u2.mem[4][8] ),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07623_ (.I(_02621_),
    .Z(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07624_ (.I(_02623_),
    .Z(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07625_ (.A1(\u2.mem[6][8] ),
    .A2(_03094_),
    .B1(_03095_),
    .B2(\u2.mem[47][8] ),
    .ZN(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07626_ (.A1(_03087_),
    .A2(_03090_),
    .A3(_03093_),
    .A4(_03096_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07627_ (.A1(_03064_),
    .A2(_03075_),
    .A3(_03086_),
    .A4(_03097_),
    .ZN(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07628_ (.A1(_01954_),
    .A2(_03013_),
    .B1(_03053_),
    .B2(_03098_),
    .ZN(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07629_ (.I(_02443_),
    .Z(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07630_ (.I(_02447_),
    .Z(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07631_ (.A1(\u2.mem[45][9] ),
    .A2(_03099_),
    .B1(_03100_),
    .B2(\u2.mem[34][9] ),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07632_ (.A1(\u2.mem[32][9] ),
    .A2(_03015_),
    .B1(_03016_),
    .B2(\u2.mem[2][9] ),
    .ZN(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07633_ (.A1(\u2.mem[40][9] ),
    .A2(_03018_),
    .B1(_03019_),
    .B2(\u2.mem[30][9] ),
    .ZN(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07634_ (.A1(\u2.mem[27][9] ),
    .A2(_03021_),
    .B1(_03022_),
    .B2(\u2.mem[35][9] ),
    .ZN(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07635_ (.A1(_03101_),
    .A2(_03102_),
    .A3(_03103_),
    .A4(_03104_),
    .ZN(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07636_ (.A1(\u2.mem[15][9] ),
    .A2(_03025_),
    .B1(_03026_),
    .B2(\u2.mem[13][9] ),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07637_ (.A1(\u2.mem[1][9] ),
    .A2(_03028_),
    .B1(_03029_),
    .B2(\u2.mem[7][9] ),
    .ZN(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07638_ (.A1(\u2.mem[16][9] ),
    .A2(_03031_),
    .B1(_03032_),
    .B2(\u2.mem[33][9] ),
    .ZN(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07639_ (.A1(\u2.mem[3][9] ),
    .A2(_03034_),
    .B(_02978_),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07640_ (.A1(_03106_),
    .A2(_03107_),
    .A3(_03108_),
    .A4(_03109_),
    .ZN(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07641_ (.I(_02502_),
    .Z(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07642_ (.I(_02504_),
    .Z(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07643_ (.A1(\u2.mem[50][9] ),
    .A2(_03111_),
    .B1(_03112_),
    .B2(\u2.mem[51][9] ),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07644_ (.I(_02508_),
    .Z(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07645_ (.I(_02510_),
    .Z(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07646_ (.A1(\u2.mem[54][9] ),
    .A2(_03114_),
    .B1(_03115_),
    .B2(\u2.mem[55][9] ),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07647_ (.A1(\u2.mem[53][9] ),
    .A2(_03039_),
    .B1(_03040_),
    .B2(\u2.mem[56][9] ),
    .ZN(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07648_ (.A1(\u2.mem[58][9] ),
    .A2(_03042_),
    .B1(_03043_),
    .B2(\u2.mem[36][9] ),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07649_ (.A1(_03113_),
    .A2(_03116_),
    .A3(_03117_),
    .A4(_03118_),
    .ZN(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07650_ (.I(_02520_),
    .Z(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07651_ (.I(_02522_),
    .Z(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07652_ (.A1(\u2.mem[44][9] ),
    .A2(_03120_),
    .B1(_03121_),
    .B2(\u2.mem[42][9] ),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07653_ (.I(_02525_),
    .Z(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07654_ (.I(_02527_),
    .Z(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07655_ (.A1(\u2.mem[14][9] ),
    .A2(_03123_),
    .B1(_03124_),
    .B2(\u2.mem[12][9] ),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07656_ (.I(_02530_),
    .Z(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07657_ (.I(_02532_),
    .Z(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07658_ (.A1(\u2.mem[49][9] ),
    .A2(_03126_),
    .B1(_03127_),
    .B2(\u2.mem[46][9] ),
    .ZN(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07659_ (.A1(\u2.mem[43][9] ),
    .A2(_03049_),
    .B1(_03050_),
    .B2(\u2.mem[20][9] ),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07660_ (.A1(_03122_),
    .A2(_03125_),
    .A3(_03128_),
    .A4(_03129_),
    .ZN(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07661_ (.A1(_03105_),
    .A2(_03110_),
    .A3(_03119_),
    .A4(_03130_),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07662_ (.I(_02558_),
    .Z(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07663_ (.I(_02560_),
    .Z(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07664_ (.A1(\u2.mem[61][9] ),
    .A2(_03132_),
    .B1(_03133_),
    .B2(\u2.mem[63][9] ),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07665_ (.A1(\u2.mem[60][9] ),
    .A2(_03055_),
    .B1(_03056_),
    .B2(\u2.mem[62][9] ),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07666_ (.A1(\u2.mem[37][9] ),
    .A2(_03058_),
    .B1(_03059_),
    .B2(\u2.mem[59][9] ),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07667_ (.A1(\u2.mem[57][9] ),
    .A2(_03061_),
    .B1(_03062_),
    .B2(\u2.mem[41][9] ),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07668_ (.A1(_03134_),
    .A2(_03135_),
    .A3(_03136_),
    .A4(_03137_),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07669_ (.I(_02572_),
    .Z(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07670_ (.I(_02574_),
    .Z(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07671_ (.A1(\u2.mem[26][9] ),
    .A2(_03139_),
    .B1(_03140_),
    .B2(\u2.mem[10][9] ),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07672_ (.A1(\u2.mem[29][9] ),
    .A2(_03066_),
    .B1(_03067_),
    .B2(\u2.mem[11][9] ),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07673_ (.A1(\u2.mem[9][9] ),
    .A2(_03069_),
    .B1(_03070_),
    .B2(\u2.mem[25][9] ),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07674_ (.A1(\u2.mem[28][9] ),
    .A2(_03072_),
    .B1(_03073_),
    .B2(\u2.mem[31][9] ),
    .ZN(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07675_ (.A1(_03141_),
    .A2(_03142_),
    .A3(_03143_),
    .A4(_03144_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07676_ (.I(_02595_),
    .Z(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07677_ (.I(_02597_),
    .Z(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07678_ (.A1(\u2.mem[23][9] ),
    .A2(_03146_),
    .B1(_03147_),
    .B2(\u2.mem[22][9] ),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07679_ (.A1(\u2.mem[17][9] ),
    .A2(_03077_),
    .B1(_03078_),
    .B2(\u2.mem[24][9] ),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07680_ (.A1(\u2.mem[52][9] ),
    .A2(_03080_),
    .B1(_03081_),
    .B2(\u2.mem[21][9] ),
    .ZN(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07681_ (.A1(\u2.mem[18][9] ),
    .A2(_03083_),
    .B1(_03084_),
    .B2(\u2.mem[19][9] ),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07682_ (.A1(_03148_),
    .A2(_03149_),
    .A3(_03150_),
    .A4(_03151_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07683_ (.I(_02626_),
    .Z(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07684_ (.I(_02628_),
    .Z(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07685_ (.A1(\u2.mem[5][9] ),
    .A2(_03153_),
    .B1(_03154_),
    .B2(\u2.mem[38][9] ),
    .ZN(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07686_ (.A1(\u2.mem[39][9] ),
    .A2(_03088_),
    .B1(_03089_),
    .B2(\u2.mem[48][9] ),
    .ZN(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07687_ (.A1(\u2.mem[8][9] ),
    .A2(_03091_),
    .B1(_03092_),
    .B2(\u2.mem[4][9] ),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07688_ (.A1(\u2.mem[6][9] ),
    .A2(_03094_),
    .B1(_03095_),
    .B2(\u2.mem[47][9] ),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07689_ (.A1(_03155_),
    .A2(_03156_),
    .A3(_03157_),
    .A4(_03158_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07690_ (.A1(_03138_),
    .A2(_03145_),
    .A3(_03152_),
    .A4(_03159_),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07691_ (.A1(_01958_),
    .A2(_03013_),
    .B1(_03131_),
    .B2(_03160_),
    .ZN(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07692_ (.A1(\u2.mem[45][10] ),
    .A2(_03099_),
    .B1(_03100_),
    .B2(\u2.mem[34][10] ),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07693_ (.A1(\u2.mem[32][10] ),
    .A2(_03015_),
    .B1(_03016_),
    .B2(\u2.mem[2][10] ),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07694_ (.A1(\u2.mem[40][10] ),
    .A2(_03018_),
    .B1(_03019_),
    .B2(\u2.mem[30][10] ),
    .ZN(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07695_ (.A1(\u2.mem[27][10] ),
    .A2(_03021_),
    .B1(_03022_),
    .B2(\u2.mem[35][10] ),
    .ZN(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07696_ (.A1(_03161_),
    .A2(_03162_),
    .A3(_03163_),
    .A4(_03164_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07697_ (.A1(\u2.mem[15][10] ),
    .A2(_03025_),
    .B1(_03026_),
    .B2(\u2.mem[13][10] ),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07698_ (.A1(\u2.mem[1][10] ),
    .A2(_03028_),
    .B1(_03029_),
    .B2(\u2.mem[7][10] ),
    .ZN(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07699_ (.A1(\u2.mem[16][10] ),
    .A2(_03031_),
    .B1(_03032_),
    .B2(\u2.mem[33][10] ),
    .ZN(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07700_ (.A1(\u2.mem[3][10] ),
    .A2(_03034_),
    .B(_02978_),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07701_ (.A1(_03166_),
    .A2(_03167_),
    .A3(_03168_),
    .A4(_03169_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07702_ (.A1(\u2.mem[50][10] ),
    .A2(_03111_),
    .B1(_03112_),
    .B2(\u2.mem[51][10] ),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07703_ (.A1(\u2.mem[54][10] ),
    .A2(_03114_),
    .B1(_03115_),
    .B2(\u2.mem[55][10] ),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07704_ (.A1(\u2.mem[53][10] ),
    .A2(_03039_),
    .B1(_03040_),
    .B2(\u2.mem[56][10] ),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07705_ (.A1(\u2.mem[58][10] ),
    .A2(_03042_),
    .B1(_03043_),
    .B2(\u2.mem[36][10] ),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07706_ (.A1(_03171_),
    .A2(_03172_),
    .A3(_03173_),
    .A4(_03174_),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07707_ (.A1(\u2.mem[44][10] ),
    .A2(_03120_),
    .B1(_03121_),
    .B2(\u2.mem[42][10] ),
    .ZN(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07708_ (.A1(\u2.mem[14][10] ),
    .A2(_03123_),
    .B1(_03124_),
    .B2(\u2.mem[12][10] ),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07709_ (.A1(\u2.mem[49][10] ),
    .A2(_03126_),
    .B1(_03127_),
    .B2(\u2.mem[46][10] ),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07710_ (.A1(\u2.mem[43][10] ),
    .A2(_03049_),
    .B1(_03050_),
    .B2(\u2.mem[20][10] ),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07711_ (.A1(_03176_),
    .A2(_03177_),
    .A3(_03178_),
    .A4(_03179_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07712_ (.A1(_03165_),
    .A2(_03170_),
    .A3(_03175_),
    .A4(_03180_),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07713_ (.A1(\u2.mem[61][10] ),
    .A2(_03132_),
    .B1(_03133_),
    .B2(\u2.mem[63][10] ),
    .ZN(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07714_ (.A1(\u2.mem[60][10] ),
    .A2(_03055_),
    .B1(_03056_),
    .B2(\u2.mem[62][10] ),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07715_ (.A1(\u2.mem[37][10] ),
    .A2(_03058_),
    .B1(_03059_),
    .B2(\u2.mem[59][10] ),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07716_ (.A1(\u2.mem[57][10] ),
    .A2(_03061_),
    .B1(_03062_),
    .B2(\u2.mem[41][10] ),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07717_ (.A1(_03182_),
    .A2(_03183_),
    .A3(_03184_),
    .A4(_03185_),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07718_ (.A1(\u2.mem[26][10] ),
    .A2(_03139_),
    .B1(_03140_),
    .B2(\u2.mem[10][10] ),
    .ZN(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07719_ (.A1(\u2.mem[29][10] ),
    .A2(_03066_),
    .B1(_03067_),
    .B2(\u2.mem[11][10] ),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07720_ (.A1(\u2.mem[9][10] ),
    .A2(_03069_),
    .B1(_03070_),
    .B2(\u2.mem[25][10] ),
    .ZN(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07721_ (.A1(\u2.mem[28][10] ),
    .A2(_03072_),
    .B1(_03073_),
    .B2(\u2.mem[31][10] ),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07722_ (.A1(_03187_),
    .A2(_03188_),
    .A3(_03189_),
    .A4(_03190_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07723_ (.A1(\u2.mem[23][10] ),
    .A2(_03146_),
    .B1(_03147_),
    .B2(\u2.mem[22][10] ),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07724_ (.A1(\u2.mem[17][10] ),
    .A2(_03077_),
    .B1(_03078_),
    .B2(\u2.mem[24][10] ),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07725_ (.A1(\u2.mem[52][10] ),
    .A2(_03080_),
    .B1(_03081_),
    .B2(\u2.mem[21][10] ),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07726_ (.A1(\u2.mem[18][10] ),
    .A2(_03083_),
    .B1(_03084_),
    .B2(\u2.mem[19][10] ),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07727_ (.A1(_03192_),
    .A2(_03193_),
    .A3(_03194_),
    .A4(_03195_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07728_ (.A1(\u2.mem[5][10] ),
    .A2(_03153_),
    .B1(_03154_),
    .B2(\u2.mem[38][10] ),
    .ZN(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07729_ (.A1(\u2.mem[39][10] ),
    .A2(_03088_),
    .B1(_03089_),
    .B2(\u2.mem[48][10] ),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07730_ (.A1(\u2.mem[8][10] ),
    .A2(_03091_),
    .B1(_03092_),
    .B2(\u2.mem[4][10] ),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07731_ (.A1(\u2.mem[6][10] ),
    .A2(_03094_),
    .B1(_03095_),
    .B2(\u2.mem[47][10] ),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07732_ (.A1(_03197_),
    .A2(_03198_),
    .A3(_03199_),
    .A4(_03200_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07733_ (.A1(_03186_),
    .A2(_03191_),
    .A3(_03196_),
    .A4(_03201_),
    .ZN(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07734_ (.A1(_01962_),
    .A2(_03013_),
    .B1(_03181_),
    .B2(_03202_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07735_ (.A1(\u2.mem[45][11] ),
    .A2(_03099_),
    .B1(_03100_),
    .B2(\u2.mem[34][11] ),
    .ZN(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07736_ (.A1(\u2.mem[32][11] ),
    .A2(_03015_),
    .B1(_03016_),
    .B2(\u2.mem[2][11] ),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07737_ (.A1(\u2.mem[40][11] ),
    .A2(_03018_),
    .B1(_03019_),
    .B2(\u2.mem[30][11] ),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07738_ (.A1(\u2.mem[27][11] ),
    .A2(_03021_),
    .B1(_03022_),
    .B2(\u2.mem[35][11] ),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07739_ (.A1(_03203_),
    .A2(_03204_),
    .A3(_03205_),
    .A4(_03206_),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07740_ (.A1(\u2.mem[15][11] ),
    .A2(_03025_),
    .B1(_03026_),
    .B2(\u2.mem[13][11] ),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07741_ (.A1(\u2.mem[1][11] ),
    .A2(_03028_),
    .B1(_03029_),
    .B2(\u2.mem[7][11] ),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07742_ (.A1(\u2.mem[16][11] ),
    .A2(_03031_),
    .B1(_03032_),
    .B2(\u2.mem[33][11] ),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07743_ (.I(_02357_),
    .Z(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07744_ (.A1(\u2.mem[3][11] ),
    .A2(_03034_),
    .B(_03211_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07745_ (.A1(_03208_),
    .A2(_03209_),
    .A3(_03210_),
    .A4(_03212_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07746_ (.A1(\u2.mem[50][11] ),
    .A2(_03111_),
    .B1(_03112_),
    .B2(\u2.mem[51][11] ),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07747_ (.A1(\u2.mem[54][11] ),
    .A2(_03114_),
    .B1(_03115_),
    .B2(\u2.mem[55][11] ),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07748_ (.A1(\u2.mem[53][11] ),
    .A2(_03039_),
    .B1(_03040_),
    .B2(\u2.mem[56][11] ),
    .ZN(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07749_ (.A1(\u2.mem[58][11] ),
    .A2(_03042_),
    .B1(_03043_),
    .B2(\u2.mem[36][11] ),
    .ZN(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07750_ (.A1(_03214_),
    .A2(_03215_),
    .A3(_03216_),
    .A4(_03217_),
    .ZN(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07751_ (.A1(\u2.mem[44][11] ),
    .A2(_03120_),
    .B1(_03121_),
    .B2(\u2.mem[42][11] ),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07752_ (.A1(\u2.mem[14][11] ),
    .A2(_03123_),
    .B1(_03124_),
    .B2(\u2.mem[12][11] ),
    .ZN(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07753_ (.A1(\u2.mem[49][11] ),
    .A2(_03126_),
    .B1(_03127_),
    .B2(\u2.mem[46][11] ),
    .ZN(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07754_ (.A1(\u2.mem[43][11] ),
    .A2(_03049_),
    .B1(_03050_),
    .B2(\u2.mem[20][11] ),
    .ZN(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07755_ (.A1(_03219_),
    .A2(_03220_),
    .A3(_03221_),
    .A4(_03222_),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07756_ (.A1(_03207_),
    .A2(_03213_),
    .A3(_03218_),
    .A4(_03223_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07757_ (.A1(\u2.mem[61][11] ),
    .A2(_03132_),
    .B1(_03133_),
    .B2(\u2.mem[63][11] ),
    .ZN(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07758_ (.A1(\u2.mem[60][11] ),
    .A2(_03055_),
    .B1(_03056_),
    .B2(\u2.mem[62][11] ),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07759_ (.A1(\u2.mem[37][11] ),
    .A2(_03058_),
    .B1(_03059_),
    .B2(\u2.mem[59][11] ),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07760_ (.A1(\u2.mem[57][11] ),
    .A2(_03061_),
    .B1(_03062_),
    .B2(\u2.mem[41][11] ),
    .ZN(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07761_ (.A1(_03225_),
    .A2(_03226_),
    .A3(_03227_),
    .A4(_03228_),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07762_ (.A1(\u2.mem[26][11] ),
    .A2(_03139_),
    .B1(_03140_),
    .B2(\u2.mem[10][11] ),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07763_ (.A1(\u2.mem[29][11] ),
    .A2(_03066_),
    .B1(_03067_),
    .B2(\u2.mem[11][11] ),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07764_ (.A1(\u2.mem[9][11] ),
    .A2(_03069_),
    .B1(_03070_),
    .B2(\u2.mem[25][11] ),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07765_ (.A1(\u2.mem[28][11] ),
    .A2(_03072_),
    .B1(_03073_),
    .B2(\u2.mem[31][11] ),
    .ZN(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07766_ (.A1(_03230_),
    .A2(_03231_),
    .A3(_03232_),
    .A4(_03233_),
    .ZN(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07767_ (.A1(\u2.mem[23][11] ),
    .A2(_03146_),
    .B1(_03147_),
    .B2(\u2.mem[22][11] ),
    .ZN(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07768_ (.A1(\u2.mem[17][11] ),
    .A2(_03077_),
    .B1(_03078_),
    .B2(\u2.mem[24][11] ),
    .ZN(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07769_ (.A1(\u2.mem[52][11] ),
    .A2(_03080_),
    .B1(_03081_),
    .B2(\u2.mem[21][11] ),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07770_ (.A1(\u2.mem[18][11] ),
    .A2(_03083_),
    .B1(_03084_),
    .B2(\u2.mem[19][11] ),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07771_ (.A1(_03235_),
    .A2(_03236_),
    .A3(_03237_),
    .A4(_03238_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07772_ (.A1(\u2.mem[5][11] ),
    .A2(_03153_),
    .B1(_03154_),
    .B2(\u2.mem[38][11] ),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07773_ (.A1(\u2.mem[39][11] ),
    .A2(_03088_),
    .B1(_03089_),
    .B2(\u2.mem[48][11] ),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07774_ (.A1(\u2.mem[8][11] ),
    .A2(_03091_),
    .B1(_03092_),
    .B2(\u2.mem[4][11] ),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07775_ (.A1(\u2.mem[6][11] ),
    .A2(_03094_),
    .B1(_03095_),
    .B2(\u2.mem[47][11] ),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07776_ (.A1(_03240_),
    .A2(_03241_),
    .A3(_03242_),
    .A4(_03243_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07777_ (.A1(_03229_),
    .A2(_03234_),
    .A3(_03239_),
    .A4(_03244_),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07778_ (.A1(_01966_),
    .A2(_03013_),
    .B1(_03224_),
    .B2(_03245_),
    .ZN(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07779_ (.I(_02360_),
    .Z(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07780_ (.A1(\u2.mem[45][12] ),
    .A2(_03099_),
    .B1(_03100_),
    .B2(\u2.mem[34][12] ),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07781_ (.I(_02385_),
    .Z(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07782_ (.I(_02395_),
    .Z(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07783_ (.A1(\u2.mem[32][12] ),
    .A2(_03248_),
    .B1(_03249_),
    .B2(\u2.mem[2][12] ),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07784_ (.I(_02405_),
    .Z(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07785_ (.I(_02414_),
    .Z(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07786_ (.A1(\u2.mem[40][12] ),
    .A2(_03251_),
    .B1(_03252_),
    .B2(\u2.mem[30][12] ),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07787_ (.I(_02427_),
    .Z(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07788_ (.I(_02435_),
    .Z(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07789_ (.A1(\u2.mem[27][12] ),
    .A2(_03254_),
    .B1(_03255_),
    .B2(\u2.mem[35][12] ),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07790_ (.A1(_03247_),
    .A2(_03250_),
    .A3(_03253_),
    .A4(_03256_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07791_ (.I(_02456_),
    .Z(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07792_ (.I(_02460_),
    .Z(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07793_ (.A1(\u2.mem[15][12] ),
    .A2(_03258_),
    .B1(_03259_),
    .B2(\u2.mem[13][12] ),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07794_ (.I(_02464_),
    .Z(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07795_ (.I(_02470_),
    .Z(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07796_ (.A1(\u2.mem[1][12] ),
    .A2(_03261_),
    .B1(_03262_),
    .B2(\u2.mem[7][12] ),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07797_ (.I(_02474_),
    .Z(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07798_ (.I(_02476_),
    .Z(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07799_ (.A1(\u2.mem[16][12] ),
    .A2(_03264_),
    .B1(_03265_),
    .B2(\u2.mem[33][12] ),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07800_ (.I(_02479_),
    .Z(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07801_ (.A1(\u2.mem[3][12] ),
    .A2(_03267_),
    .B(_03211_),
    .ZN(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07802_ (.A1(_03260_),
    .A2(_03263_),
    .A3(_03266_),
    .A4(_03268_),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07803_ (.A1(\u2.mem[50][12] ),
    .A2(_03111_),
    .B1(_03112_),
    .B2(\u2.mem[51][12] ),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07804_ (.A1(\u2.mem[54][12] ),
    .A2(_03114_),
    .B1(_03115_),
    .B2(\u2.mem[55][12] ),
    .ZN(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07805_ (.I(_02485_),
    .Z(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07806_ (.I(_02488_),
    .Z(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07807_ (.A1(\u2.mem[53][12] ),
    .A2(_03272_),
    .B1(_03273_),
    .B2(\u2.mem[56][12] ),
    .ZN(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07808_ (.I(_02494_),
    .Z(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07809_ (.I(_02499_),
    .Z(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07810_ (.A1(\u2.mem[58][12] ),
    .A2(_03275_),
    .B1(_03276_),
    .B2(\u2.mem[36][12] ),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07811_ (.A1(_03270_),
    .A2(_03271_),
    .A3(_03274_),
    .A4(_03277_),
    .ZN(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07812_ (.A1(\u2.mem[44][12] ),
    .A2(_03120_),
    .B1(_03121_),
    .B2(\u2.mem[42][12] ),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07813_ (.A1(\u2.mem[14][12] ),
    .A2(_03123_),
    .B1(_03124_),
    .B2(\u2.mem[12][12] ),
    .ZN(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07814_ (.A1(\u2.mem[49][12] ),
    .A2(_03126_),
    .B1(_03127_),
    .B2(\u2.mem[46][12] ),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07815_ (.I(_02514_),
    .Z(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07816_ (.I(_02516_),
    .Z(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07817_ (.A1(\u2.mem[43][12] ),
    .A2(_03282_),
    .B1(_03283_),
    .B2(\u2.mem[20][12] ),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07818_ (.A1(_03279_),
    .A2(_03280_),
    .A3(_03281_),
    .A4(_03284_),
    .ZN(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07819_ (.A1(_03257_),
    .A2(_03269_),
    .A3(_03278_),
    .A4(_03285_),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07820_ (.A1(\u2.mem[61][12] ),
    .A2(_03132_),
    .B1(_03133_),
    .B2(\u2.mem[63][12] ),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07821_ (.I(_02545_),
    .Z(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07822_ (.I(_02548_),
    .Z(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07823_ (.A1(\u2.mem[60][12] ),
    .A2(_03288_),
    .B1(_03289_),
    .B2(\u2.mem[62][12] ),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07824_ (.I(_02539_),
    .Z(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07825_ (.I(_02541_),
    .Z(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07826_ (.A1(\u2.mem[37][12] ),
    .A2(_03291_),
    .B1(_03292_),
    .B2(\u2.mem[59][12] ),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07827_ (.I(_02553_),
    .Z(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07828_ (.I(_02555_),
    .Z(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07829_ (.A1(\u2.mem[57][12] ),
    .A2(_03294_),
    .B1(_03295_),
    .B2(\u2.mem[41][12] ),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07830_ (.A1(_03287_),
    .A2(_03290_),
    .A3(_03293_),
    .A4(_03296_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07831_ (.A1(\u2.mem[26][12] ),
    .A2(_03139_),
    .B1(_03140_),
    .B2(\u2.mem[10][12] ),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07832_ (.I(_02564_),
    .Z(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07833_ (.I(_02569_),
    .Z(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07834_ (.A1(\u2.mem[29][12] ),
    .A2(_03299_),
    .B1(_03300_),
    .B2(\u2.mem[11][12] ),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07835_ (.I(_02579_),
    .Z(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07836_ (.I(_02581_),
    .Z(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07837_ (.A1(\u2.mem[9][12] ),
    .A2(_03302_),
    .B1(_03303_),
    .B2(\u2.mem[25][12] ),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07838_ (.I(_02584_),
    .Z(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07839_ (.I(_02586_),
    .Z(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07840_ (.A1(\u2.mem[28][12] ),
    .A2(_03305_),
    .B1(_03306_),
    .B2(\u2.mem[31][12] ),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07841_ (.A1(_03298_),
    .A2(_03301_),
    .A3(_03304_),
    .A4(_03307_),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07842_ (.A1(\u2.mem[23][12] ),
    .A2(_03146_),
    .B1(_03147_),
    .B2(\u2.mem[22][12] ),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07843_ (.I(_02590_),
    .Z(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07844_ (.I(_02592_),
    .Z(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07845_ (.A1(\u2.mem[17][12] ),
    .A2(_03310_),
    .B1(_03311_),
    .B2(\u2.mem[24][12] ),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07846_ (.I(_02600_),
    .Z(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07847_ (.I(_02602_),
    .Z(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07848_ (.A1(\u2.mem[52][12] ),
    .A2(_03313_),
    .B1(_03314_),
    .B2(\u2.mem[21][12] ),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07849_ (.I(_02605_),
    .Z(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07850_ (.I(_02607_),
    .Z(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07851_ (.A1(\u2.mem[18][12] ),
    .A2(_03316_),
    .B1(_03317_),
    .B2(\u2.mem[19][12] ),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07852_ (.A1(_03309_),
    .A2(_03312_),
    .A3(_03315_),
    .A4(_03318_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07853_ (.A1(\u2.mem[5][12] ),
    .A2(_03153_),
    .B1(_03154_),
    .B2(\u2.mem[38][12] ),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07854_ (.I(_02616_),
    .Z(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07855_ (.I(_02618_),
    .Z(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07856_ (.A1(\u2.mem[39][12] ),
    .A2(_03321_),
    .B1(_03322_),
    .B2(\u2.mem[48][12] ),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07857_ (.I(_02611_),
    .Z(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07858_ (.I(_02613_),
    .Z(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07859_ (.A1(\u2.mem[8][12] ),
    .A2(_03324_),
    .B1(_03325_),
    .B2(\u2.mem[4][12] ),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07860_ (.I(_02621_),
    .Z(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07861_ (.I(_02623_),
    .Z(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07862_ (.A1(\u2.mem[6][12] ),
    .A2(_03327_),
    .B1(_03328_),
    .B2(\u2.mem[47][12] ),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07863_ (.A1(_03320_),
    .A2(_03323_),
    .A3(_03326_),
    .A4(_03329_),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07864_ (.A1(_03297_),
    .A2(_03308_),
    .A3(_03319_),
    .A4(_03330_),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07865_ (.A1(_01969_),
    .A2(_03246_),
    .B1(_03286_),
    .B2(_03331_),
    .ZN(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07866_ (.A1(\u2.mem[45][13] ),
    .A2(_02444_),
    .B1(_02448_),
    .B2(\u2.mem[34][13] ),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07867_ (.A1(\u2.mem[32][13] ),
    .A2(_03248_),
    .B1(_03249_),
    .B2(\u2.mem[2][13] ),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07868_ (.A1(\u2.mem[40][13] ),
    .A2(_03251_),
    .B1(_03252_),
    .B2(\u2.mem[30][13] ),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07869_ (.A1(\u2.mem[27][13] ),
    .A2(_03254_),
    .B1(_03255_),
    .B2(\u2.mem[35][13] ),
    .ZN(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07870_ (.A1(_03332_),
    .A2(_03333_),
    .A3(_03334_),
    .A4(_03335_),
    .ZN(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07871_ (.A1(\u2.mem[15][13] ),
    .A2(_03258_),
    .B1(_03259_),
    .B2(\u2.mem[13][13] ),
    .ZN(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07872_ (.A1(\u2.mem[1][13] ),
    .A2(_03261_),
    .B1(_03262_),
    .B2(\u2.mem[7][13] ),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07873_ (.A1(\u2.mem[16][13] ),
    .A2(_03264_),
    .B1(_03265_),
    .B2(\u2.mem[33][13] ),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07874_ (.A1(\u2.mem[3][13] ),
    .A2(_03267_),
    .B(_03211_),
    .ZN(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07875_ (.A1(_03337_),
    .A2(_03338_),
    .A3(_03339_),
    .A4(_03340_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07876_ (.A1(\u2.mem[50][13] ),
    .A2(_02503_),
    .B1(_02505_),
    .B2(\u2.mem[51][13] ),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07877_ (.A1(\u2.mem[54][13] ),
    .A2(_02509_),
    .B1(_02511_),
    .B2(\u2.mem[55][13] ),
    .ZN(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07878_ (.A1(\u2.mem[53][13] ),
    .A2(_03272_),
    .B1(_03273_),
    .B2(\u2.mem[56][13] ),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07879_ (.A1(\u2.mem[58][13] ),
    .A2(_03275_),
    .B1(_03276_),
    .B2(\u2.mem[36][13] ),
    .ZN(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07880_ (.A1(_03342_),
    .A2(_03343_),
    .A3(_03344_),
    .A4(_03345_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07881_ (.A1(\u2.mem[44][13] ),
    .A2(_02521_),
    .B1(_02523_),
    .B2(\u2.mem[42][13] ),
    .ZN(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07882_ (.A1(\u2.mem[14][13] ),
    .A2(_02526_),
    .B1(_02528_),
    .B2(\u2.mem[12][13] ),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07883_ (.A1(\u2.mem[49][13] ),
    .A2(_02531_),
    .B1(_02533_),
    .B2(\u2.mem[46][13] ),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07884_ (.A1(\u2.mem[43][13] ),
    .A2(_03282_),
    .B1(_03283_),
    .B2(\u2.mem[20][13] ),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07885_ (.A1(_03347_),
    .A2(_03348_),
    .A3(_03349_),
    .A4(_03350_),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07886_ (.A1(_03336_),
    .A2(_03341_),
    .A3(_03346_),
    .A4(_03351_),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07887_ (.A1(\u2.mem[61][13] ),
    .A2(_02559_),
    .B1(_02561_),
    .B2(\u2.mem[63][13] ),
    .ZN(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07888_ (.A1(\u2.mem[60][13] ),
    .A2(_03288_),
    .B1(_03289_),
    .B2(\u2.mem[62][13] ),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07889_ (.A1(\u2.mem[37][13] ),
    .A2(_03291_),
    .B1(_03292_),
    .B2(\u2.mem[59][13] ),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07890_ (.A1(\u2.mem[57][13] ),
    .A2(_03294_),
    .B1(_03295_),
    .B2(\u2.mem[41][13] ),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07891_ (.A1(_03353_),
    .A2(_03354_),
    .A3(_03355_),
    .A4(_03356_),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07892_ (.A1(\u2.mem[26][13] ),
    .A2(_02573_),
    .B1(_02575_),
    .B2(\u2.mem[10][13] ),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07893_ (.A1(\u2.mem[29][13] ),
    .A2(_03299_),
    .B1(_03300_),
    .B2(\u2.mem[11][13] ),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07894_ (.A1(\u2.mem[9][13] ),
    .A2(_03302_),
    .B1(_03303_),
    .B2(\u2.mem[25][13] ),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07895_ (.A1(\u2.mem[28][13] ),
    .A2(_03305_),
    .B1(_03306_),
    .B2(\u2.mem[31][13] ),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07896_ (.A1(_03358_),
    .A2(_03359_),
    .A3(_03360_),
    .A4(_03361_),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07897_ (.A1(\u2.mem[23][13] ),
    .A2(_02596_),
    .B1(_02598_),
    .B2(\u2.mem[22][13] ),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07898_ (.A1(\u2.mem[17][13] ),
    .A2(_03310_),
    .B1(_03311_),
    .B2(\u2.mem[24][13] ),
    .ZN(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07899_ (.A1(\u2.mem[52][13] ),
    .A2(_03313_),
    .B1(_03314_),
    .B2(\u2.mem[21][13] ),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07900_ (.A1(\u2.mem[18][13] ),
    .A2(_03316_),
    .B1(_03317_),
    .B2(\u2.mem[19][13] ),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07901_ (.A1(_03363_),
    .A2(_03364_),
    .A3(_03365_),
    .A4(_03366_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07902_ (.A1(\u2.mem[5][13] ),
    .A2(_02627_),
    .B1(_02629_),
    .B2(\u2.mem[38][13] ),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07903_ (.A1(\u2.mem[39][13] ),
    .A2(_03321_),
    .B1(_03322_),
    .B2(\u2.mem[48][13] ),
    .ZN(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07904_ (.A1(\u2.mem[8][13] ),
    .A2(_03324_),
    .B1(_03325_),
    .B2(\u2.mem[4][13] ),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07905_ (.A1(\u2.mem[6][13] ),
    .A2(_03327_),
    .B1(_03328_),
    .B2(\u2.mem[47][13] ),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07906_ (.A1(_03368_),
    .A2(_03369_),
    .A3(_03370_),
    .A4(_03371_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07907_ (.A1(_03357_),
    .A2(_03362_),
    .A3(_03367_),
    .A4(_03372_),
    .ZN(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07908_ (.A1(_01973_),
    .A2(_03246_),
    .B1(_03352_),
    .B2(_03373_),
    .ZN(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07909_ (.A1(\u2.mem[45][14] ),
    .A2(_02444_),
    .B1(_02448_),
    .B2(\u2.mem[34][14] ),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07910_ (.A1(\u2.mem[32][14] ),
    .A2(_03248_),
    .B1(_03249_),
    .B2(\u2.mem[2][14] ),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07911_ (.A1(\u2.mem[40][14] ),
    .A2(_03251_),
    .B1(_03252_),
    .B2(\u2.mem[30][14] ),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07912_ (.A1(\u2.mem[27][14] ),
    .A2(_03254_),
    .B1(_03255_),
    .B2(\u2.mem[35][14] ),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07913_ (.A1(_03374_),
    .A2(_03375_),
    .A3(_03376_),
    .A4(_03377_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07914_ (.A1(\u2.mem[15][14] ),
    .A2(_03258_),
    .B1(_03259_),
    .B2(\u2.mem[13][14] ),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07915_ (.A1(\u2.mem[1][14] ),
    .A2(_03261_),
    .B1(_03262_),
    .B2(\u2.mem[7][14] ),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07916_ (.A1(\u2.mem[16][14] ),
    .A2(_03264_),
    .B1(_03265_),
    .B2(\u2.mem[33][14] ),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07917_ (.A1(\u2.mem[3][14] ),
    .A2(_03267_),
    .B(_03211_),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07918_ (.A1(_03379_),
    .A2(_03380_),
    .A3(_03381_),
    .A4(_03382_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07919_ (.A1(\u2.mem[50][14] ),
    .A2(_02503_),
    .B1(_02505_),
    .B2(\u2.mem[51][14] ),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07920_ (.A1(\u2.mem[54][14] ),
    .A2(_02509_),
    .B1(_02511_),
    .B2(\u2.mem[55][14] ),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07921_ (.A1(\u2.mem[53][14] ),
    .A2(_03272_),
    .B1(_03273_),
    .B2(\u2.mem[56][14] ),
    .ZN(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07922_ (.A1(\u2.mem[58][14] ),
    .A2(_03275_),
    .B1(_03276_),
    .B2(\u2.mem[36][14] ),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07923_ (.A1(_03384_),
    .A2(_03385_),
    .A3(_03386_),
    .A4(_03387_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07924_ (.A1(\u2.mem[44][14] ),
    .A2(_02521_),
    .B1(_02523_),
    .B2(\u2.mem[42][14] ),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07925_ (.A1(\u2.mem[14][14] ),
    .A2(_02526_),
    .B1(_02528_),
    .B2(\u2.mem[12][14] ),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07926_ (.A1(\u2.mem[49][14] ),
    .A2(_02531_),
    .B1(_02533_),
    .B2(\u2.mem[46][14] ),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07927_ (.A1(\u2.mem[43][14] ),
    .A2(_03282_),
    .B1(_03283_),
    .B2(\u2.mem[20][14] ),
    .ZN(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07928_ (.A1(_03389_),
    .A2(_03390_),
    .A3(_03391_),
    .A4(_03392_),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07929_ (.A1(_03378_),
    .A2(_03383_),
    .A3(_03388_),
    .A4(_03393_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07930_ (.A1(\u2.mem[61][14] ),
    .A2(_02559_),
    .B1(_02561_),
    .B2(\u2.mem[63][14] ),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07931_ (.A1(\u2.mem[60][14] ),
    .A2(_03288_),
    .B1(_03289_),
    .B2(\u2.mem[62][14] ),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07932_ (.A1(\u2.mem[37][14] ),
    .A2(_03291_),
    .B1(_03292_),
    .B2(\u2.mem[59][14] ),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07933_ (.A1(\u2.mem[57][14] ),
    .A2(_03294_),
    .B1(_03295_),
    .B2(\u2.mem[41][14] ),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07934_ (.A1(_03395_),
    .A2(_03396_),
    .A3(_03397_),
    .A4(_03398_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07935_ (.A1(\u2.mem[26][14] ),
    .A2(_02573_),
    .B1(_02575_),
    .B2(\u2.mem[10][14] ),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07936_ (.A1(\u2.mem[29][14] ),
    .A2(_03299_),
    .B1(_03300_),
    .B2(\u2.mem[11][14] ),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07937_ (.A1(\u2.mem[9][14] ),
    .A2(_03302_),
    .B1(_03303_),
    .B2(\u2.mem[25][14] ),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07938_ (.A1(\u2.mem[28][14] ),
    .A2(_03305_),
    .B1(_03306_),
    .B2(\u2.mem[31][14] ),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07939_ (.A1(_03400_),
    .A2(_03401_),
    .A3(_03402_),
    .A4(_03403_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07940_ (.A1(\u2.mem[23][14] ),
    .A2(_02596_),
    .B1(_02598_),
    .B2(\u2.mem[22][14] ),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07941_ (.A1(\u2.mem[17][14] ),
    .A2(_03310_),
    .B1(_03311_),
    .B2(\u2.mem[24][14] ),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07942_ (.A1(\u2.mem[52][14] ),
    .A2(_03313_),
    .B1(_03314_),
    .B2(\u2.mem[21][14] ),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07943_ (.A1(\u2.mem[18][14] ),
    .A2(_03316_),
    .B1(_03317_),
    .B2(\u2.mem[19][14] ),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07944_ (.A1(_03405_),
    .A2(_03406_),
    .A3(_03407_),
    .A4(_03408_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07945_ (.A1(\u2.mem[5][14] ),
    .A2(_02627_),
    .B1(_02629_),
    .B2(\u2.mem[38][14] ),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07946_ (.A1(\u2.mem[39][14] ),
    .A2(_03321_),
    .B1(_03322_),
    .B2(\u2.mem[48][14] ),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07947_ (.A1(\u2.mem[8][14] ),
    .A2(_03324_),
    .B1(_03325_),
    .B2(\u2.mem[4][14] ),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07948_ (.A1(\u2.mem[6][14] ),
    .A2(_03327_),
    .B1(_03328_),
    .B2(\u2.mem[47][14] ),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07949_ (.A1(_03410_),
    .A2(_03411_),
    .A3(_03412_),
    .A4(_03413_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07950_ (.A1(_03399_),
    .A2(_03404_),
    .A3(_03409_),
    .A4(_03414_),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07951_ (.A1(_01976_),
    .A2(_03246_),
    .B1(_03394_),
    .B2(_03415_),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07952_ (.A1(\u2.mem[45][15] ),
    .A2(_02444_),
    .B1(_02448_),
    .B2(\u2.mem[34][15] ),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07953_ (.A1(\u2.mem[32][15] ),
    .A2(_03248_),
    .B1(_03249_),
    .B2(\u2.mem[2][15] ),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07954_ (.A1(\u2.mem[40][15] ),
    .A2(_03251_),
    .B1(_03252_),
    .B2(\u2.mem[30][15] ),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07955_ (.A1(\u2.mem[27][15] ),
    .A2(_03254_),
    .B1(_03255_),
    .B2(\u2.mem[35][15] ),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07956_ (.A1(_03416_),
    .A2(_03417_),
    .A3(_03418_),
    .A4(_03419_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07957_ (.A1(\u2.mem[15][15] ),
    .A2(_03258_),
    .B1(_03259_),
    .B2(\u2.mem[13][15] ),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07958_ (.A1(\u2.mem[1][15] ),
    .A2(_03261_),
    .B1(_03262_),
    .B2(\u2.mem[7][15] ),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07959_ (.A1(\u2.mem[16][15] ),
    .A2(_03264_),
    .B1(_03265_),
    .B2(\u2.mem[33][15] ),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07960_ (.A1(\u2.mem[3][15] ),
    .A2(_03267_),
    .B(_02358_),
    .ZN(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07961_ (.A1(_03421_),
    .A2(_03422_),
    .A3(_03423_),
    .A4(_03424_),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07962_ (.A1(\u2.mem[50][15] ),
    .A2(_02503_),
    .B1(_02505_),
    .B2(\u2.mem[51][15] ),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07963_ (.A1(\u2.mem[54][15] ),
    .A2(_02509_),
    .B1(_02511_),
    .B2(\u2.mem[55][15] ),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07964_ (.A1(\u2.mem[53][15] ),
    .A2(_03272_),
    .B1(_03273_),
    .B2(\u2.mem[56][15] ),
    .ZN(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07965_ (.A1(\u2.mem[58][15] ),
    .A2(_03275_),
    .B1(_03276_),
    .B2(\u2.mem[36][15] ),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07966_ (.A1(_03426_),
    .A2(_03427_),
    .A3(_03428_),
    .A4(_03429_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07967_ (.A1(\u2.mem[44][15] ),
    .A2(_02521_),
    .B1(_02523_),
    .B2(\u2.mem[42][15] ),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07968_ (.A1(\u2.mem[14][15] ),
    .A2(_02526_),
    .B1(_02528_),
    .B2(\u2.mem[12][15] ),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07969_ (.A1(\u2.mem[49][15] ),
    .A2(_02531_),
    .B1(_02533_),
    .B2(\u2.mem[46][15] ),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07970_ (.A1(\u2.mem[43][15] ),
    .A2(_03282_),
    .B1(_03283_),
    .B2(\u2.mem[20][15] ),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07971_ (.A1(_03431_),
    .A2(_03432_),
    .A3(_03433_),
    .A4(_03434_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07972_ (.A1(_03420_),
    .A2(_03425_),
    .A3(_03430_),
    .A4(_03435_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07973_ (.A1(\u2.mem[61][15] ),
    .A2(_02559_),
    .B1(_02561_),
    .B2(\u2.mem[63][15] ),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07974_ (.A1(\u2.mem[60][15] ),
    .A2(_03288_),
    .B1(_03289_),
    .B2(\u2.mem[62][15] ),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07975_ (.A1(\u2.mem[37][15] ),
    .A2(_03291_),
    .B1(_03292_),
    .B2(\u2.mem[59][15] ),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07976_ (.A1(\u2.mem[57][15] ),
    .A2(_03294_),
    .B1(_03295_),
    .B2(\u2.mem[41][15] ),
    .ZN(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07977_ (.A1(_03437_),
    .A2(_03438_),
    .A3(_03439_),
    .A4(_03440_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07978_ (.A1(\u2.mem[26][15] ),
    .A2(_02573_),
    .B1(_02575_),
    .B2(\u2.mem[10][15] ),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07979_ (.A1(\u2.mem[29][15] ),
    .A2(_03299_),
    .B1(_03300_),
    .B2(\u2.mem[11][15] ),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07980_ (.A1(\u2.mem[9][15] ),
    .A2(_03302_),
    .B1(_03303_),
    .B2(\u2.mem[25][15] ),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07981_ (.A1(\u2.mem[28][15] ),
    .A2(_03305_),
    .B1(_03306_),
    .B2(\u2.mem[31][15] ),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07982_ (.A1(_03442_),
    .A2(_03443_),
    .A3(_03444_),
    .A4(_03445_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07983_ (.A1(\u2.mem[23][15] ),
    .A2(_02596_),
    .B1(_02598_),
    .B2(\u2.mem[22][15] ),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07984_ (.A1(\u2.mem[17][15] ),
    .A2(_03310_),
    .B1(_03311_),
    .B2(\u2.mem[24][15] ),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07985_ (.A1(\u2.mem[52][15] ),
    .A2(_03313_),
    .B1(_03314_),
    .B2(\u2.mem[21][15] ),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07986_ (.A1(\u2.mem[18][15] ),
    .A2(_03316_),
    .B1(_03317_),
    .B2(\u2.mem[19][15] ),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07987_ (.A1(_03447_),
    .A2(_03448_),
    .A3(_03449_),
    .A4(_03450_),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07988_ (.A1(\u2.mem[5][15] ),
    .A2(_02627_),
    .B1(_02629_),
    .B2(\u2.mem[38][15] ),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07989_ (.A1(\u2.mem[39][15] ),
    .A2(_03321_),
    .B1(_03322_),
    .B2(\u2.mem[48][15] ),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07990_ (.A1(\u2.mem[8][15] ),
    .A2(_03324_),
    .B1(_03325_),
    .B2(\u2.mem[4][15] ),
    .ZN(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07991_ (.A1(\u2.mem[6][15] ),
    .A2(_03327_),
    .B1(_03328_),
    .B2(\u2.mem[47][15] ),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07992_ (.A1(_03452_),
    .A2(_03453_),
    .A3(_03454_),
    .A4(_03455_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07993_ (.A1(_03441_),
    .A2(_03446_),
    .A3(_03451_),
    .A4(_03456_),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07994_ (.A1(_01980_),
    .A2(_03246_),
    .B1(_03436_),
    .B2(_03457_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07995_ (.A1(_01562_),
    .A2(_01575_),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07996_ (.I(_01613_),
    .Z(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07997_ (.A1(\u2.active_mem[4] ),
    .A2(_03458_),
    .B1(_03459_),
    .B2(\u2.active_mem[5] ),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07998_ (.I(_01547_),
    .Z(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07999_ (.I(_01665_),
    .Z(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08000_ (.A1(\u2.active_mem[7] ),
    .A2(_03461_),
    .B1(_03462_),
    .B2(\u2.active_mem[6] ),
    .ZN(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08001_ (.A1(_03460_),
    .A2(_03463_),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08002_ (.A1(\u2.active_mem[11] ),
    .A2(_03461_),
    .B1(_03462_),
    .B2(\u2.active_mem[10] ),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08003_ (.A1(\u2.active_mem[8] ),
    .A2(_03458_),
    .B1(_03459_),
    .B2(\u2.active_mem[9] ),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08004_ (.A1(_03465_),
    .A2(_03466_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08005_ (.A1(_01591_),
    .A2(_03464_),
    .B1(_03467_),
    .B2(_01678_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08006_ (.A1(\u2.active_mem[12] ),
    .A2(_03458_),
    .B1(_03459_),
    .B2(\u2.active_mem[13] ),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08007_ (.A1(\u2.active_mem[15] ),
    .A2(_03461_),
    .B1(_03462_),
    .B2(\u2.active_mem[14] ),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08008_ (.A1(_03469_),
    .A2(_03470_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08009_ (.A1(\u2.active_mem[3] ),
    .A2(_03461_),
    .B1(_03462_),
    .B2(\u2.active_mem[2] ),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08010_ (.A1(\u2.active_mem[0] ),
    .A2(_03458_),
    .B1(_03459_),
    .B2(\u2.active_mem[1] ),
    .ZN(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08011_ (.A1(_03472_),
    .A2(_03473_),
    .B(_01549_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08012_ (.A1(_01612_),
    .A2(_03471_),
    .B(_03474_),
    .ZN(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08013_ (.A1(_03468_),
    .A2(_03475_),
    .ZN(_05992_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08014_ (.I(\u3.enable ),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08015_ (.A1(\u3.data ),
    .A2(_03476_),
    .ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08016_ (.I(\mem_address_trans[4].data_sync ),
    .Z(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08017_ (.I(\mem_address_trans[6].data_sync ),
    .Z(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _08018_ (.A1(_03477_),
    .A2(\mem_address_trans[5].data_sync ),
    .A3(_03478_),
    .A4(\mem_address_trans[7].data_sync ),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08019_ (.I(_03479_),
    .Z(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08020_ (.I(\mem_address_trans[1].data_sync ),
    .Z(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08021_ (.I(\mem_address_trans[0].data_sync ),
    .Z(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08022_ (.A1(\mem_address_trans[2].data_sync ),
    .A2(\mem_address_trans[3].data_sync ),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08023_ (.A1(\mem_write_n_trans.data_sync ),
    .A2(\mem_address_trans[9].data_sync ),
    .A3(\mem_address_trans[8].data_sync ),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08024_ (.A1(_03483_),
    .A2(_03484_),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08025_ (.A1(_03481_),
    .A2(_03482_),
    .A3(_03485_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08026_ (.I(_03486_),
    .Z(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08027_ (.A1(_03480_),
    .A2(_03487_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08028_ (.I(_03488_),
    .Z(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08029_ (.I(_03489_),
    .Z(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08030_ (.I(\data_in_trans[0].data_sync ),
    .Z(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08031_ (.I(_03491_),
    .Z(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08032_ (.I(_03488_),
    .Z(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08033_ (.I(_03493_),
    .Z(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08034_ (.A1(_03492_),
    .A2(_03494_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08035_ (.A1(_01545_),
    .A2(_03490_),
    .B(_03495_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08036_ (.I(\data_in_trans[1].data_sync ),
    .Z(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08037_ (.I(_03496_),
    .Z(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08038_ (.A1(_03497_),
    .A2(_03494_),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08039_ (.A1(_01727_),
    .A2(_03490_),
    .B(_03498_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08040_ (.I(\data_in_trans[2].data_sync ),
    .Z(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08041_ (.I(_03499_),
    .Z(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08042_ (.A1(_03500_),
    .A2(_03494_),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08043_ (.A1(_01769_),
    .A2(_03490_),
    .B(_03501_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08044_ (.I(\data_in_trans[3].data_sync ),
    .Z(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08045_ (.I(_03502_),
    .Z(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08046_ (.A1(_03503_),
    .A2(_03494_),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08047_ (.A1(_01809_),
    .A2(_03490_),
    .B(_03504_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08048_ (.I(_03489_),
    .Z(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08049_ (.I(\data_in_trans[4].data_sync ),
    .Z(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08050_ (.I(_03506_),
    .Z(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08051_ (.I(_03493_),
    .Z(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08052_ (.A1(_03507_),
    .A2(_03508_),
    .ZN(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08053_ (.A1(_01844_),
    .A2(_03505_),
    .B(_03509_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08054_ (.I(\data_in_trans[5].data_sync ),
    .Z(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08055_ (.I(_03510_),
    .Z(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08056_ (.A1(_03511_),
    .A2(_03508_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08057_ (.A1(_01878_),
    .A2(_03505_),
    .B(_03512_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08058_ (.I(\data_in_trans[6].data_sync ),
    .Z(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08059_ (.A1(_03513_),
    .A2(_03508_),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08060_ (.A1(_01945_),
    .A2(_03505_),
    .B(_03514_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08061_ (.I(\data_in_trans[7].data_sync ),
    .Z(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08062_ (.A1(_03515_),
    .A2(_03508_),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08063_ (.A1(_01951_),
    .A2(_03505_),
    .B(_03516_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08064_ (.I(_03489_),
    .Z(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08065_ (.I(\data_in_trans[8].data_sync ),
    .Z(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08066_ (.I(_03493_),
    .Z(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08067_ (.A1(_03518_),
    .A2(_03519_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08068_ (.A1(_01954_),
    .A2(_03517_),
    .B(_03520_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08069_ (.I(\data_in_trans[9].data_sync ),
    .Z(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08070_ (.A1(_03521_),
    .A2(_03519_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08071_ (.A1(_01958_),
    .A2(_03517_),
    .B(_03522_),
    .ZN(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08072_ (.I(\data_in_trans[10].data_sync ),
    .Z(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08073_ (.A1(_03523_),
    .A2(_03519_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08074_ (.A1(_01962_),
    .A2(_03517_),
    .B(_03524_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08075_ (.I(\data_in_trans[11].data_sync ),
    .Z(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08076_ (.A1(_03525_),
    .A2(_03519_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08077_ (.A1(_01966_),
    .A2(_03517_),
    .B(_03526_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08078_ (.I(_03489_),
    .Z(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08079_ (.I(\data_in_trans[12].data_sync ),
    .Z(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08080_ (.I(_03493_),
    .Z(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08081_ (.A1(_03528_),
    .A2(_03529_),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08082_ (.A1(_01969_),
    .A2(_03527_),
    .B(_03530_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08083_ (.I(\data_in_trans[13].data_sync ),
    .Z(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08084_ (.A1(_03531_),
    .A2(_03529_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08085_ (.A1(_01973_),
    .A2(_03527_),
    .B(_03532_),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08086_ (.I(\data_in_trans[14].data_sync ),
    .Z(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08087_ (.A1(_03533_),
    .A2(_03529_),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08088_ (.A1(_01976_),
    .A2(_03527_),
    .B(_03534_),
    .ZN(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08089_ (.I(\data_in_trans[15].data_sync ),
    .Z(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08090_ (.A1(_03535_),
    .A2(_03529_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08091_ (.A1(_01980_),
    .A2(_03527_),
    .B(_03536_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08092_ (.A1(\output_active_hold[3] ),
    .A2(\output_active_hold[2] ),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08093_ (.A1(\u2.driver_enable ),
    .A2(\output_active_hold[1] ),
    .A3(\output_active_hold[0] ),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08094_ (.A1(_03537_),
    .A2(_03538_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08095_ (.I(_03492_),
    .Z(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08096_ (.I(_03484_),
    .Z(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08097_ (.A1(_03479_),
    .A2(_03540_),
    .Z(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08098_ (.I(_03541_),
    .Z(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08099_ (.I(\mem_address_trans[0].data_sync ),
    .ZN(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08100_ (.A1(_03481_),
    .A2(_03543_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08101_ (.A1(_03483_),
    .A2(_03542_),
    .A3(_03544_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08102_ (.I(_03545_),
    .Z(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08103_ (.I0(_03539_),
    .I1(\u2.mem[1][0] ),
    .S(_03546_),
    .Z(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08104_ (.I(_03547_),
    .Z(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08105_ (.I(_03497_),
    .Z(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08106_ (.I0(_03548_),
    .I1(\u2.mem[1][1] ),
    .S(_03546_),
    .Z(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08107_ (.I(_03549_),
    .Z(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08108_ (.I(_03500_),
    .Z(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08109_ (.I0(_03550_),
    .I1(\u2.mem[1][2] ),
    .S(_03546_),
    .Z(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08110_ (.I(_03551_),
    .Z(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08111_ (.I(_03503_),
    .Z(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08112_ (.I0(_03552_),
    .I1(\u2.mem[1][3] ),
    .S(_03546_),
    .Z(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08113_ (.I(_03553_),
    .Z(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08114_ (.I(_03507_),
    .Z(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08115_ (.I(_03545_),
    .Z(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08116_ (.I0(_03554_),
    .I1(\u2.mem[1][4] ),
    .S(_03555_),
    .Z(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08117_ (.I(_03556_),
    .Z(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08118_ (.I(_03511_),
    .Z(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08119_ (.I0(_03557_),
    .I1(\u2.mem[1][5] ),
    .S(_03555_),
    .Z(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08120_ (.I(_03558_),
    .Z(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08121_ (.I(_03513_),
    .Z(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08122_ (.I0(_03559_),
    .I1(\u2.mem[1][6] ),
    .S(_03555_),
    .Z(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08123_ (.I(_03560_),
    .Z(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08124_ (.I(_03515_),
    .Z(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08125_ (.I0(_03561_),
    .I1(\u2.mem[1][7] ),
    .S(_03555_),
    .Z(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08126_ (.I(_03562_),
    .Z(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08127_ (.I(_03518_),
    .Z(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08128_ (.I(_03545_),
    .Z(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08129_ (.I0(_03563_),
    .I1(\u2.mem[1][8] ),
    .S(_03564_),
    .Z(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08130_ (.I(_03565_),
    .Z(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08131_ (.I(_03521_),
    .Z(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08132_ (.I0(_03566_),
    .I1(\u2.mem[1][9] ),
    .S(_03564_),
    .Z(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08133_ (.I(_03567_),
    .Z(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08134_ (.I(_03523_),
    .Z(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08135_ (.I0(_03568_),
    .I1(\u2.mem[1][10] ),
    .S(_03564_),
    .Z(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08136_ (.I(_03569_),
    .Z(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08137_ (.I(_03525_),
    .Z(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08138_ (.I0(_03570_),
    .I1(\u2.mem[1][11] ),
    .S(_03564_),
    .Z(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08139_ (.I(_03571_),
    .Z(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08140_ (.I(_03528_),
    .Z(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08141_ (.I(_03545_),
    .Z(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08142_ (.I0(_03572_),
    .I1(\u2.mem[1][12] ),
    .S(_03573_),
    .Z(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08143_ (.I(_03574_),
    .Z(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08144_ (.I(_03531_),
    .Z(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08145_ (.I0(_03575_),
    .I1(\u2.mem[1][13] ),
    .S(_03573_),
    .Z(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08146_ (.I(_03576_),
    .Z(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08147_ (.I(_03533_),
    .Z(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08148_ (.I0(_03577_),
    .I1(\u2.mem[1][14] ),
    .S(_03573_),
    .Z(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08149_ (.I(_03578_),
    .Z(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08150_ (.I(_03535_),
    .Z(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08151_ (.I0(_03579_),
    .I1(\u2.mem[1][15] ),
    .S(_03573_),
    .Z(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08152_ (.I(_03580_),
    .Z(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08153_ (.A1(_03481_),
    .A2(_03543_),
    .ZN(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08154_ (.A1(_03485_),
    .A2(_03581_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08155_ (.I(_03582_),
    .Z(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08156_ (.A1(_03480_),
    .A2(_03583_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08157_ (.I(_03584_),
    .Z(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08158_ (.I0(_03539_),
    .I1(\u2.mem[2][0] ),
    .S(_03585_),
    .Z(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08159_ (.I(_03586_),
    .Z(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08160_ (.I0(_03548_),
    .I1(\u2.mem[2][1] ),
    .S(_03585_),
    .Z(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08161_ (.I(_03587_),
    .Z(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08162_ (.I0(_03550_),
    .I1(\u2.mem[2][2] ),
    .S(_03585_),
    .Z(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08163_ (.I(_03588_),
    .Z(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08164_ (.I0(_03552_),
    .I1(\u2.mem[2][3] ),
    .S(_03585_),
    .Z(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08165_ (.I(_03589_),
    .Z(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08166_ (.I(_03584_),
    .Z(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08167_ (.I0(_03554_),
    .I1(\u2.mem[2][4] ),
    .S(_03590_),
    .Z(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08168_ (.I(_03591_),
    .Z(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08169_ (.I0(_03557_),
    .I1(\u2.mem[2][5] ),
    .S(_03590_),
    .Z(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08170_ (.I(_03592_),
    .Z(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08171_ (.I0(_03559_),
    .I1(\u2.mem[2][6] ),
    .S(_03590_),
    .Z(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08172_ (.I(_03593_),
    .Z(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08173_ (.I0(_03561_),
    .I1(\u2.mem[2][7] ),
    .S(_03590_),
    .Z(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08174_ (.I(_03594_),
    .Z(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08175_ (.I(_03584_),
    .Z(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08176_ (.I0(_03563_),
    .I1(\u2.mem[2][8] ),
    .S(_03595_),
    .Z(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08177_ (.I(_03596_),
    .Z(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08178_ (.I0(_03566_),
    .I1(\u2.mem[2][9] ),
    .S(_03595_),
    .Z(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08179_ (.I(_03597_),
    .Z(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08180_ (.I0(_03568_),
    .I1(\u2.mem[2][10] ),
    .S(_03595_),
    .Z(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08181_ (.I(_03598_),
    .Z(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08182_ (.I0(_03570_),
    .I1(\u2.mem[2][11] ),
    .S(_03595_),
    .Z(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08183_ (.I(_03599_),
    .Z(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08184_ (.I(_03584_),
    .Z(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08185_ (.I0(_03572_),
    .I1(\u2.mem[2][12] ),
    .S(_03600_),
    .Z(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08186_ (.I(_03601_),
    .Z(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08187_ (.I0(_03575_),
    .I1(\u2.mem[2][13] ),
    .S(_03600_),
    .Z(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08188_ (.I(_03602_),
    .Z(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08189_ (.I0(_03577_),
    .I1(\u2.mem[2][14] ),
    .S(_03600_),
    .Z(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08190_ (.I(_03603_),
    .Z(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08191_ (.I0(_03579_),
    .I1(\u2.mem[2][15] ),
    .S(_03600_),
    .Z(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08192_ (.I(_03604_),
    .Z(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _08193_ (.I(\mem_address_trans[1].data_sync ),
    .Z(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _08194_ (.I(_03482_),
    .Z(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08195_ (.I(_03541_),
    .Z(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08196_ (.A1(_03605_),
    .A2(_03606_),
    .A3(_03483_),
    .A4(_03607_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08197_ (.I(_03608_),
    .Z(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08198_ (.I0(_03539_),
    .I1(\u2.mem[3][0] ),
    .S(_03609_),
    .Z(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08199_ (.I(_03610_),
    .Z(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08200_ (.I0(_03548_),
    .I1(\u2.mem[3][1] ),
    .S(_03609_),
    .Z(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08201_ (.I(_03611_),
    .Z(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08202_ (.I0(_03550_),
    .I1(\u2.mem[3][2] ),
    .S(_03609_),
    .Z(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08203_ (.I(_03612_),
    .Z(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08204_ (.I0(_03552_),
    .I1(\u2.mem[3][3] ),
    .S(_03609_),
    .Z(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08205_ (.I(_03613_),
    .Z(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08206_ (.I(_03608_),
    .Z(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08207_ (.I0(_03554_),
    .I1(\u2.mem[3][4] ),
    .S(_03614_),
    .Z(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08208_ (.I(_03615_),
    .Z(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08209_ (.I0(_03557_),
    .I1(\u2.mem[3][5] ),
    .S(_03614_),
    .Z(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08210_ (.I(_03616_),
    .Z(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08211_ (.I0(_03559_),
    .I1(\u2.mem[3][6] ),
    .S(_03614_),
    .Z(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08212_ (.I(_03617_),
    .Z(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08213_ (.I0(_03561_),
    .I1(\u2.mem[3][7] ),
    .S(_03614_),
    .Z(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08214_ (.I(_03618_),
    .Z(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08215_ (.I(_03608_),
    .Z(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08216_ (.I0(_03563_),
    .I1(\u2.mem[3][8] ),
    .S(_03619_),
    .Z(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08217_ (.I(_03620_),
    .Z(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08218_ (.I0(_03566_),
    .I1(\u2.mem[3][9] ),
    .S(_03619_),
    .Z(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08219_ (.I(_03621_),
    .Z(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08220_ (.I0(_03568_),
    .I1(\u2.mem[3][10] ),
    .S(_03619_),
    .Z(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08221_ (.I(_03622_),
    .Z(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08222_ (.I0(_03570_),
    .I1(\u2.mem[3][11] ),
    .S(_03619_),
    .Z(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08223_ (.I(_03623_),
    .Z(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08224_ (.I(_03608_),
    .Z(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08225_ (.I0(_03572_),
    .I1(\u2.mem[3][12] ),
    .S(_03624_),
    .Z(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08226_ (.I(_03625_),
    .Z(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08227_ (.I0(_03575_),
    .I1(\u2.mem[3][13] ),
    .S(_03624_),
    .Z(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08228_ (.I(_03626_),
    .Z(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08229_ (.I0(_03577_),
    .I1(\u2.mem[3][14] ),
    .S(_03624_),
    .Z(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08230_ (.I(_03627_),
    .Z(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08231_ (.I0(_03579_),
    .I1(\u2.mem[3][15] ),
    .S(_03624_),
    .Z(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08232_ (.I(_03628_),
    .Z(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08233_ (.A1(\mem_address_trans[1].data_sync ),
    .A2(\mem_address_trans[0].data_sync ),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08234_ (.I(_03629_),
    .Z(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08235_ (.I(\mem_address_trans[2].data_sync ),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08236_ (.A1(_03631_),
    .A2(\mem_address_trans[3].data_sync ),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08237_ (.I(_03632_),
    .Z(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08238_ (.A1(_03630_),
    .A2(_03542_),
    .A3(_03633_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08239_ (.I(_03634_),
    .Z(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08240_ (.I0(_03539_),
    .I1(\u2.mem[4][0] ),
    .S(_03635_),
    .Z(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08241_ (.I(_03636_),
    .Z(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08242_ (.I0(_03548_),
    .I1(\u2.mem[4][1] ),
    .S(_03635_),
    .Z(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08243_ (.I(_03637_),
    .Z(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08244_ (.I0(_03550_),
    .I1(\u2.mem[4][2] ),
    .S(_03635_),
    .Z(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08245_ (.I(_03638_),
    .Z(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08246_ (.I0(_03552_),
    .I1(\u2.mem[4][3] ),
    .S(_03635_),
    .Z(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08247_ (.I(_03639_),
    .Z(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08248_ (.I(_03634_),
    .Z(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08249_ (.I0(_03554_),
    .I1(\u2.mem[4][4] ),
    .S(_03640_),
    .Z(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08250_ (.I(_03641_),
    .Z(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08251_ (.I0(_03557_),
    .I1(\u2.mem[4][5] ),
    .S(_03640_),
    .Z(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08252_ (.I(_03642_),
    .Z(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08253_ (.I0(_03559_),
    .I1(\u2.mem[4][6] ),
    .S(_03640_),
    .Z(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08254_ (.I(_03643_),
    .Z(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08255_ (.I0(_03561_),
    .I1(\u2.mem[4][7] ),
    .S(_03640_),
    .Z(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08256_ (.I(_03644_),
    .Z(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08257_ (.I(_03634_),
    .Z(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08258_ (.I0(_03563_),
    .I1(\u2.mem[4][8] ),
    .S(_03645_),
    .Z(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08259_ (.I(_03646_),
    .Z(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08260_ (.I0(_03566_),
    .I1(\u2.mem[4][9] ),
    .S(_03645_),
    .Z(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08261_ (.I(_03647_),
    .Z(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08262_ (.I0(_03568_),
    .I1(\u2.mem[4][10] ),
    .S(_03645_),
    .Z(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08263_ (.I(_03648_),
    .Z(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08264_ (.I0(_03570_),
    .I1(\u2.mem[4][11] ),
    .S(_03645_),
    .Z(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08265_ (.I(_03649_),
    .Z(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08266_ (.I(_03634_),
    .Z(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08267_ (.I0(_03572_),
    .I1(\u2.mem[4][12] ),
    .S(_03650_),
    .Z(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08268_ (.I(_03651_),
    .Z(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08269_ (.I0(_03575_),
    .I1(\u2.mem[4][13] ),
    .S(_03650_),
    .Z(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08270_ (.I(_03652_),
    .Z(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08271_ (.I0(_03577_),
    .I1(\u2.mem[4][14] ),
    .S(_03650_),
    .Z(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08272_ (.I(_03653_),
    .Z(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08273_ (.I0(_03579_),
    .I1(\u2.mem[4][15] ),
    .S(_03650_),
    .Z(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08274_ (.I(_03654_),
    .Z(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08275_ (.I(_03491_),
    .Z(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08276_ (.I(_03655_),
    .Z(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08277_ (.I(_03656_),
    .Z(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08278_ (.I(_03541_),
    .Z(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08279_ (.A1(_03658_),
    .A2(_03544_),
    .A3(_03633_),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08280_ (.I(_03659_),
    .Z(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08281_ (.I0(_03657_),
    .I1(\u2.mem[5][0] ),
    .S(_03660_),
    .Z(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08282_ (.I(_03661_),
    .Z(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08283_ (.I(_03496_),
    .Z(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08284_ (.I(_03662_),
    .Z(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08285_ (.I(_03663_),
    .Z(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08286_ (.I0(_03664_),
    .I1(\u2.mem[5][1] ),
    .S(_03660_),
    .Z(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08287_ (.I(_03665_),
    .Z(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08288_ (.I(_03499_),
    .Z(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08289_ (.I(_03666_),
    .Z(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08290_ (.I(_03667_),
    .Z(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08291_ (.I0(_03668_),
    .I1(\u2.mem[5][2] ),
    .S(_03660_),
    .Z(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08292_ (.I(_03669_),
    .Z(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08293_ (.I(_03502_),
    .Z(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08294_ (.I(_03670_),
    .Z(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08295_ (.I(_03671_),
    .Z(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08296_ (.I0(_03672_),
    .I1(\u2.mem[5][3] ),
    .S(_03660_),
    .Z(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08297_ (.I(_03673_),
    .Z(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08298_ (.I(_03506_),
    .Z(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08299_ (.I(_03674_),
    .Z(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08300_ (.I(_03675_),
    .Z(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08301_ (.I(_03659_),
    .Z(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08302_ (.I0(_03676_),
    .I1(\u2.mem[5][4] ),
    .S(_03677_),
    .Z(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08303_ (.I(_03678_),
    .Z(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08304_ (.I(_03510_),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08305_ (.I(_03679_),
    .Z(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08306_ (.I(_03680_),
    .Z(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08307_ (.I0(_03681_),
    .I1(\u2.mem[5][5] ),
    .S(_03677_),
    .Z(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08308_ (.I(_03682_),
    .Z(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08309_ (.I(\data_in_trans[6].data_sync ),
    .Z(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08310_ (.I(_03683_),
    .Z(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08311_ (.I(_03684_),
    .Z(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08312_ (.I0(_03685_),
    .I1(\u2.mem[5][6] ),
    .S(_03677_),
    .Z(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08313_ (.I(_03686_),
    .Z(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08314_ (.I(\data_in_trans[7].data_sync ),
    .Z(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08315_ (.I(_03687_),
    .Z(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08316_ (.I(_03688_),
    .Z(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08317_ (.I0(_03689_),
    .I1(\u2.mem[5][7] ),
    .S(_03677_),
    .Z(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08318_ (.I(_03690_),
    .Z(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08319_ (.I(\data_in_trans[8].data_sync ),
    .Z(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08320_ (.I(_03691_),
    .Z(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08321_ (.I(_03692_),
    .Z(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08322_ (.I(_03659_),
    .Z(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08323_ (.I0(_03693_),
    .I1(\u2.mem[5][8] ),
    .S(_03694_),
    .Z(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08324_ (.I(_03695_),
    .Z(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08325_ (.I(\data_in_trans[9].data_sync ),
    .Z(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08326_ (.I(_03696_),
    .Z(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08327_ (.I(_03697_),
    .Z(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08328_ (.I0(_03698_),
    .I1(\u2.mem[5][9] ),
    .S(_03694_),
    .Z(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08329_ (.I(_03699_),
    .Z(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08330_ (.I(\data_in_trans[10].data_sync ),
    .Z(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08331_ (.I(_03700_),
    .Z(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08332_ (.I(_03701_),
    .Z(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08333_ (.I0(_03702_),
    .I1(\u2.mem[5][10] ),
    .S(_03694_),
    .Z(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08334_ (.I(_03703_),
    .Z(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08335_ (.I(\data_in_trans[11].data_sync ),
    .Z(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08336_ (.I(_03704_),
    .Z(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08337_ (.I(_03705_),
    .Z(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08338_ (.I0(_03706_),
    .I1(\u2.mem[5][11] ),
    .S(_03694_),
    .Z(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08339_ (.I(_03707_),
    .Z(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08340_ (.I(\data_in_trans[12].data_sync ),
    .Z(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08341_ (.I(_03708_),
    .Z(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08342_ (.I(_03709_),
    .Z(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08343_ (.I(_03659_),
    .Z(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08344_ (.I0(_03710_),
    .I1(\u2.mem[5][12] ),
    .S(_03711_),
    .Z(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08345_ (.I(_03712_),
    .Z(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08346_ (.I(\data_in_trans[13].data_sync ),
    .Z(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08347_ (.I(_03713_),
    .Z(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08348_ (.I(_03714_),
    .Z(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08349_ (.I0(_03715_),
    .I1(\u2.mem[5][13] ),
    .S(_03711_),
    .Z(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08350_ (.I(_03716_),
    .Z(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08351_ (.I(\data_in_trans[14].data_sync ),
    .Z(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08352_ (.I(_03717_),
    .Z(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08353_ (.I(_03718_),
    .Z(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08354_ (.I0(_03719_),
    .I1(\u2.mem[5][14] ),
    .S(_03711_),
    .Z(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08355_ (.I(_03720_),
    .Z(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08356_ (.I(\data_in_trans[15].data_sync ),
    .Z(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08357_ (.I(_03721_),
    .Z(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08358_ (.I(_03722_),
    .Z(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08359_ (.I0(_03723_),
    .I1(\u2.mem[5][15] ),
    .S(_03711_),
    .Z(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08360_ (.I(_03724_),
    .Z(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08361_ (.I(_03481_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08362_ (.A1(_03725_),
    .A2(_03606_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08363_ (.A1(_03658_),
    .A2(_03726_),
    .A3(_03633_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08364_ (.I(_03727_),
    .Z(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08365_ (.I0(_03657_),
    .I1(\u2.mem[6][0] ),
    .S(_03728_),
    .Z(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08366_ (.I(_03729_),
    .Z(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08367_ (.I0(_03664_),
    .I1(\u2.mem[6][1] ),
    .S(_03728_),
    .Z(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08368_ (.I(_03730_),
    .Z(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08369_ (.I0(_03668_),
    .I1(\u2.mem[6][2] ),
    .S(_03728_),
    .Z(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08370_ (.I(_03731_),
    .Z(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08371_ (.I0(_03672_),
    .I1(\u2.mem[6][3] ),
    .S(_03728_),
    .Z(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08372_ (.I(_03732_),
    .Z(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08373_ (.I(_03727_),
    .Z(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08374_ (.I0(_03676_),
    .I1(\u2.mem[6][4] ),
    .S(_03733_),
    .Z(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08375_ (.I(_03734_),
    .Z(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08376_ (.I0(_03681_),
    .I1(\u2.mem[6][5] ),
    .S(_03733_),
    .Z(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08377_ (.I(_03735_),
    .Z(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08378_ (.I0(_03685_),
    .I1(\u2.mem[6][6] ),
    .S(_03733_),
    .Z(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08379_ (.I(_03736_),
    .Z(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08380_ (.I0(_03689_),
    .I1(\u2.mem[6][7] ),
    .S(_03733_),
    .Z(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08381_ (.I(_03737_),
    .Z(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08382_ (.I(_03727_),
    .Z(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08383_ (.I0(_03693_),
    .I1(\u2.mem[6][8] ),
    .S(_03738_),
    .Z(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08384_ (.I(_03739_),
    .Z(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08385_ (.I0(_03698_),
    .I1(\u2.mem[6][9] ),
    .S(_03738_),
    .Z(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08386_ (.I(_03740_),
    .Z(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08387_ (.I0(_03702_),
    .I1(\u2.mem[6][10] ),
    .S(_03738_),
    .Z(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08388_ (.I(_03741_),
    .Z(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08389_ (.I0(_03706_),
    .I1(\u2.mem[6][11] ),
    .S(_03738_),
    .Z(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08390_ (.I(_03742_),
    .Z(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08391_ (.I(_03727_),
    .Z(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08392_ (.I0(_03710_),
    .I1(\u2.mem[6][12] ),
    .S(_03743_),
    .Z(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08393_ (.I(_03744_),
    .Z(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08394_ (.I0(_03715_),
    .I1(\u2.mem[6][13] ),
    .S(_03743_),
    .Z(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08395_ (.I(_03745_),
    .Z(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08396_ (.I0(_03719_),
    .I1(\u2.mem[6][14] ),
    .S(_03743_),
    .Z(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08397_ (.I(_03746_),
    .Z(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08398_ (.I0(_03723_),
    .I1(\u2.mem[6][15] ),
    .S(_03743_),
    .Z(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08399_ (.I(_03747_),
    .Z(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08400_ (.A1(_03605_),
    .A2(_03482_),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08401_ (.I(_03484_),
    .Z(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08402_ (.A1(_03749_),
    .A2(_03632_),
    .ZN(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08403_ (.A1(_03748_),
    .A2(_03750_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08404_ (.I(_03751_),
    .Z(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08405_ (.A1(_03480_),
    .A2(_03752_),
    .ZN(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08406_ (.I(_03753_),
    .Z(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08407_ (.I0(_03657_),
    .I1(\u2.mem[7][0] ),
    .S(_03754_),
    .Z(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08408_ (.I(_03755_),
    .Z(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08409_ (.I0(_03664_),
    .I1(\u2.mem[7][1] ),
    .S(_03754_),
    .Z(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08410_ (.I(_03756_),
    .Z(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08411_ (.I0(_03668_),
    .I1(\u2.mem[7][2] ),
    .S(_03754_),
    .Z(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08412_ (.I(_03757_),
    .Z(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08413_ (.I0(_03672_),
    .I1(\u2.mem[7][3] ),
    .S(_03754_),
    .Z(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08414_ (.I(_03758_),
    .Z(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08415_ (.I(_03753_),
    .Z(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08416_ (.I0(_03676_),
    .I1(\u2.mem[7][4] ),
    .S(_03759_),
    .Z(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08417_ (.I(_03760_),
    .Z(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08418_ (.I0(_03681_),
    .I1(\u2.mem[7][5] ),
    .S(_03759_),
    .Z(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08419_ (.I(_03761_),
    .Z(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08420_ (.I0(_03685_),
    .I1(\u2.mem[7][6] ),
    .S(_03759_),
    .Z(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08421_ (.I(_03762_),
    .Z(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08422_ (.I0(_03689_),
    .I1(\u2.mem[7][7] ),
    .S(_03759_),
    .Z(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08423_ (.I(_03763_),
    .Z(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08424_ (.I(_03753_),
    .Z(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08425_ (.I0(_03693_),
    .I1(\u2.mem[7][8] ),
    .S(_03764_),
    .Z(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08426_ (.I(_03765_),
    .Z(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08427_ (.I0(_03698_),
    .I1(\u2.mem[7][9] ),
    .S(_03764_),
    .Z(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08428_ (.I(_03766_),
    .Z(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08429_ (.I0(_03702_),
    .I1(\u2.mem[7][10] ),
    .S(_03764_),
    .Z(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08430_ (.I(_03767_),
    .Z(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08431_ (.I0(_03706_),
    .I1(\u2.mem[7][11] ),
    .S(_03764_),
    .Z(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08432_ (.I(_03768_),
    .Z(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08433_ (.I(_03753_),
    .Z(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08434_ (.I0(_03710_),
    .I1(\u2.mem[7][12] ),
    .S(_03769_),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08435_ (.I(_03770_),
    .Z(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08436_ (.I0(_03715_),
    .I1(\u2.mem[7][13] ),
    .S(_03769_),
    .Z(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08437_ (.I(_03771_),
    .Z(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08438_ (.I0(_03719_),
    .I1(\u2.mem[7][14] ),
    .S(_03769_),
    .Z(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08439_ (.I(_03772_),
    .Z(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08440_ (.I0(_03723_),
    .I1(\u2.mem[7][15] ),
    .S(_03769_),
    .Z(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08441_ (.I(_03773_),
    .Z(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08442_ (.I(\mem_address_trans[3].data_sync ),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08443_ (.A1(\mem_address_trans[2].data_sync ),
    .A2(_03774_),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08444_ (.I(_03775_),
    .Z(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08445_ (.A1(_03630_),
    .A2(_03542_),
    .A3(_03776_),
    .ZN(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08446_ (.I(_03777_),
    .Z(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08447_ (.I0(_03657_),
    .I1(\u2.mem[8][0] ),
    .S(_03778_),
    .Z(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08448_ (.I(_03779_),
    .Z(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08449_ (.I0(_03664_),
    .I1(\u2.mem[8][1] ),
    .S(_03778_),
    .Z(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08450_ (.I(_03780_),
    .Z(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08451_ (.I0(_03668_),
    .I1(\u2.mem[8][2] ),
    .S(_03778_),
    .Z(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08452_ (.I(_03781_),
    .Z(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08453_ (.I0(_03672_),
    .I1(\u2.mem[8][3] ),
    .S(_03778_),
    .Z(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08454_ (.I(_03782_),
    .Z(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08455_ (.I(_03777_),
    .Z(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08456_ (.I0(_03676_),
    .I1(\u2.mem[8][4] ),
    .S(_03783_),
    .Z(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08457_ (.I(_03784_),
    .Z(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08458_ (.I0(_03681_),
    .I1(\u2.mem[8][5] ),
    .S(_03783_),
    .Z(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08459_ (.I(_03785_),
    .Z(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08460_ (.I0(_03685_),
    .I1(\u2.mem[8][6] ),
    .S(_03783_),
    .Z(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08461_ (.I(_03786_),
    .Z(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08462_ (.I0(_03689_),
    .I1(\u2.mem[8][7] ),
    .S(_03783_),
    .Z(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08463_ (.I(_03787_),
    .Z(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08464_ (.I(_03777_),
    .Z(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08465_ (.I0(_03693_),
    .I1(\u2.mem[8][8] ),
    .S(_03788_),
    .Z(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08466_ (.I(_03789_),
    .Z(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08467_ (.I0(_03698_),
    .I1(\u2.mem[8][9] ),
    .S(_03788_),
    .Z(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08468_ (.I(_03790_),
    .Z(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08469_ (.I0(_03702_),
    .I1(\u2.mem[8][10] ),
    .S(_03788_),
    .Z(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08470_ (.I(_03791_),
    .Z(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08471_ (.I0(_03706_),
    .I1(\u2.mem[8][11] ),
    .S(_03788_),
    .Z(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08472_ (.I(_03792_),
    .Z(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08473_ (.I(_03777_),
    .Z(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08474_ (.I0(_03710_),
    .I1(\u2.mem[8][12] ),
    .S(_03793_),
    .Z(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08475_ (.I(_03794_),
    .Z(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08476_ (.I0(_03715_),
    .I1(\u2.mem[8][13] ),
    .S(_03793_),
    .Z(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08477_ (.I(_03795_),
    .Z(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08478_ (.I0(_03719_),
    .I1(\u2.mem[8][14] ),
    .S(_03793_),
    .Z(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08479_ (.I(_03796_),
    .Z(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08480_ (.I0(_03723_),
    .I1(\u2.mem[8][15] ),
    .S(_03793_),
    .Z(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08481_ (.I(_03797_),
    .Z(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08482_ (.I(_03656_),
    .Z(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08483_ (.A1(_03658_),
    .A2(_03544_),
    .A3(_03776_),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08484_ (.I(_03799_),
    .Z(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08485_ (.I0(_03798_),
    .I1(\u2.mem[9][0] ),
    .S(_03800_),
    .Z(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08486_ (.I(_03801_),
    .Z(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08487_ (.I(_03663_),
    .Z(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08488_ (.I0(_03802_),
    .I1(\u2.mem[9][1] ),
    .S(_03800_),
    .Z(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08489_ (.I(_03803_),
    .Z(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08490_ (.I(_03667_),
    .Z(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08491_ (.I0(_03804_),
    .I1(\u2.mem[9][2] ),
    .S(_03800_),
    .Z(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08492_ (.I(_03805_),
    .Z(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08493_ (.I(_03671_),
    .Z(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08494_ (.I0(_03806_),
    .I1(\u2.mem[9][3] ),
    .S(_03800_),
    .Z(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08495_ (.I(_03807_),
    .Z(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08496_ (.I(_03675_),
    .Z(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08497_ (.I(_03799_),
    .Z(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08498_ (.I0(_03808_),
    .I1(\u2.mem[9][4] ),
    .S(_03809_),
    .Z(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08499_ (.I(_03810_),
    .Z(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08500_ (.I(_03680_),
    .Z(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08501_ (.I0(_03811_),
    .I1(\u2.mem[9][5] ),
    .S(_03809_),
    .Z(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08502_ (.I(_03812_),
    .Z(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08503_ (.I(_03684_),
    .Z(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08504_ (.I0(_03813_),
    .I1(\u2.mem[9][6] ),
    .S(_03809_),
    .Z(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08505_ (.I(_03814_),
    .Z(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08506_ (.I(_03688_),
    .Z(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08507_ (.I0(_03815_),
    .I1(\u2.mem[9][7] ),
    .S(_03809_),
    .Z(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08508_ (.I(_03816_),
    .Z(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08509_ (.I(_03692_),
    .Z(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08510_ (.I(_03799_),
    .Z(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08511_ (.I0(_03817_),
    .I1(\u2.mem[9][8] ),
    .S(_03818_),
    .Z(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08512_ (.I(_03819_),
    .Z(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08513_ (.I(_03697_),
    .Z(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08514_ (.I0(_03820_),
    .I1(\u2.mem[9][9] ),
    .S(_03818_),
    .Z(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08515_ (.I(_03821_),
    .Z(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08516_ (.I(_03701_),
    .Z(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08517_ (.I0(_03822_),
    .I1(\u2.mem[9][10] ),
    .S(_03818_),
    .Z(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08518_ (.I(_03823_),
    .Z(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08519_ (.I(_03705_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08520_ (.I0(_03824_),
    .I1(\u2.mem[9][11] ),
    .S(_03818_),
    .Z(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08521_ (.I(_03825_),
    .Z(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08522_ (.I(_03709_),
    .Z(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08523_ (.I(_03799_),
    .Z(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08524_ (.I0(_03826_),
    .I1(\u2.mem[9][12] ),
    .S(_03827_),
    .Z(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08525_ (.I(_03828_),
    .Z(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08526_ (.I(_03714_),
    .Z(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08527_ (.I0(_03829_),
    .I1(\u2.mem[9][13] ),
    .S(_03827_),
    .Z(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08528_ (.I(_03830_),
    .Z(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08529_ (.I(_03718_),
    .Z(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08530_ (.I0(_03831_),
    .I1(\u2.mem[9][14] ),
    .S(_03827_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08531_ (.I(_03832_),
    .Z(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08532_ (.I(_03722_),
    .Z(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08533_ (.I0(_03833_),
    .I1(\u2.mem[9][15] ),
    .S(_03827_),
    .Z(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08534_ (.I(_03834_),
    .Z(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08535_ (.A1(_03658_),
    .A2(_03726_),
    .A3(_03776_),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08536_ (.I(_03835_),
    .Z(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08537_ (.I0(_03798_),
    .I1(\u2.mem[10][0] ),
    .S(_03836_),
    .Z(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08538_ (.I(_03837_),
    .Z(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08539_ (.I0(_03802_),
    .I1(\u2.mem[10][1] ),
    .S(_03836_),
    .Z(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08540_ (.I(_03838_),
    .Z(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08541_ (.I0(_03804_),
    .I1(\u2.mem[10][2] ),
    .S(_03836_),
    .Z(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08542_ (.I(_03839_),
    .Z(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08543_ (.I0(_03806_),
    .I1(\u2.mem[10][3] ),
    .S(_03836_),
    .Z(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08544_ (.I(_03840_),
    .Z(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08545_ (.I(_03835_),
    .Z(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08546_ (.I0(_03808_),
    .I1(\u2.mem[10][4] ),
    .S(_03841_),
    .Z(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08547_ (.I(_03842_),
    .Z(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08548_ (.I0(_03811_),
    .I1(\u2.mem[10][5] ),
    .S(_03841_),
    .Z(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08549_ (.I(_03843_),
    .Z(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08550_ (.I0(_03813_),
    .I1(\u2.mem[10][6] ),
    .S(_03841_),
    .Z(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08551_ (.I(_03844_),
    .Z(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08552_ (.I0(_03815_),
    .I1(\u2.mem[10][7] ),
    .S(_03841_),
    .Z(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08553_ (.I(_03845_),
    .Z(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08554_ (.I(_03835_),
    .Z(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08555_ (.I0(_03817_),
    .I1(\u2.mem[10][8] ),
    .S(_03846_),
    .Z(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08556_ (.I(_03847_),
    .Z(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08557_ (.I0(_03820_),
    .I1(\u2.mem[10][9] ),
    .S(_03846_),
    .Z(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08558_ (.I(_03848_),
    .Z(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08559_ (.I0(_03822_),
    .I1(\u2.mem[10][10] ),
    .S(_03846_),
    .Z(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08560_ (.I(_03849_),
    .Z(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08561_ (.I0(_03824_),
    .I1(\u2.mem[10][11] ),
    .S(_03846_),
    .Z(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08562_ (.I(_03850_),
    .Z(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08563_ (.I(_03835_),
    .Z(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08564_ (.I0(_03826_),
    .I1(\u2.mem[10][12] ),
    .S(_03851_),
    .Z(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08565_ (.I(_03852_),
    .Z(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08566_ (.I0(_03829_),
    .I1(\u2.mem[10][13] ),
    .S(_03851_),
    .Z(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08567_ (.I(_03853_),
    .Z(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08568_ (.I0(_03831_),
    .I1(\u2.mem[10][14] ),
    .S(_03851_),
    .Z(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08569_ (.I(_03854_),
    .Z(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08570_ (.I0(_03833_),
    .I1(\u2.mem[10][15] ),
    .S(_03851_),
    .Z(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08571_ (.I(_03855_),
    .Z(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08572_ (.A1(_03605_),
    .A2(_03606_),
    .A3(_03607_),
    .A4(_03776_),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08573_ (.I(_03856_),
    .Z(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08574_ (.I0(_03798_),
    .I1(\u2.mem[11][0] ),
    .S(_03857_),
    .Z(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08575_ (.I(_03858_),
    .Z(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08576_ (.I0(_03802_),
    .I1(\u2.mem[11][1] ),
    .S(_03857_),
    .Z(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08577_ (.I(_03859_),
    .Z(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08578_ (.I0(_03804_),
    .I1(\u2.mem[11][2] ),
    .S(_03857_),
    .Z(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08579_ (.I(_03860_),
    .Z(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08580_ (.I0(_03806_),
    .I1(\u2.mem[11][3] ),
    .S(_03857_),
    .Z(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08581_ (.I(_03861_),
    .Z(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08582_ (.I(_03856_),
    .Z(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08583_ (.I0(_03808_),
    .I1(\u2.mem[11][4] ),
    .S(_03862_),
    .Z(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08584_ (.I(_03863_),
    .Z(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08585_ (.I0(_03811_),
    .I1(\u2.mem[11][5] ),
    .S(_03862_),
    .Z(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08586_ (.I(_03864_),
    .Z(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08587_ (.I0(_03813_),
    .I1(\u2.mem[11][6] ),
    .S(_03862_),
    .Z(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08588_ (.I(_03865_),
    .Z(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08589_ (.I0(_03815_),
    .I1(\u2.mem[11][7] ),
    .S(_03862_),
    .Z(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08590_ (.I(_03866_),
    .Z(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08591_ (.I(_03856_),
    .Z(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08592_ (.I0(_03817_),
    .I1(\u2.mem[11][8] ),
    .S(_03867_),
    .Z(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08593_ (.I(_03868_),
    .Z(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08594_ (.I0(_03820_),
    .I1(\u2.mem[11][9] ),
    .S(_03867_),
    .Z(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08595_ (.I(_03869_),
    .Z(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08596_ (.I0(_03822_),
    .I1(\u2.mem[11][10] ),
    .S(_03867_),
    .Z(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08597_ (.I(_03870_),
    .Z(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08598_ (.I0(_03824_),
    .I1(\u2.mem[11][11] ),
    .S(_03867_),
    .Z(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08599_ (.I(_03871_),
    .Z(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08600_ (.I(_03856_),
    .Z(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08601_ (.I0(_03826_),
    .I1(\u2.mem[11][12] ),
    .S(_03872_),
    .Z(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08602_ (.I(_03873_),
    .Z(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08603_ (.I0(_03829_),
    .I1(\u2.mem[11][13] ),
    .S(_03872_),
    .Z(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08604_ (.I(_03874_),
    .Z(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08605_ (.I0(_03831_),
    .I1(\u2.mem[11][14] ),
    .S(_03872_),
    .Z(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08606_ (.I(_03875_),
    .Z(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08607_ (.I0(_03833_),
    .I1(\u2.mem[11][15] ),
    .S(_03872_),
    .Z(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08608_ (.I(_03876_),
    .Z(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08609_ (.A1(_03631_),
    .A2(_03774_),
    .ZN(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08610_ (.I(_03877_),
    .Z(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08611_ (.A1(_03630_),
    .A2(_03542_),
    .A3(_03878_),
    .ZN(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08612_ (.I(_03879_),
    .Z(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08613_ (.I0(_03798_),
    .I1(\u2.mem[12][0] ),
    .S(_03880_),
    .Z(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08614_ (.I(_03881_),
    .Z(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08615_ (.I0(_03802_),
    .I1(\u2.mem[12][1] ),
    .S(_03880_),
    .Z(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08616_ (.I(_03882_),
    .Z(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08617_ (.I0(_03804_),
    .I1(\u2.mem[12][2] ),
    .S(_03880_),
    .Z(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08618_ (.I(_03883_),
    .Z(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08619_ (.I0(_03806_),
    .I1(\u2.mem[12][3] ),
    .S(_03880_),
    .Z(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08620_ (.I(_03884_),
    .Z(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08621_ (.I(_03879_),
    .Z(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08622_ (.I0(_03808_),
    .I1(\u2.mem[12][4] ),
    .S(_03885_),
    .Z(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08623_ (.I(_03886_),
    .Z(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08624_ (.I0(_03811_),
    .I1(\u2.mem[12][5] ),
    .S(_03885_),
    .Z(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08625_ (.I(_03887_),
    .Z(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08626_ (.I0(_03813_),
    .I1(\u2.mem[12][6] ),
    .S(_03885_),
    .Z(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08627_ (.I(_03888_),
    .Z(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08628_ (.I0(_03815_),
    .I1(\u2.mem[12][7] ),
    .S(_03885_),
    .Z(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08629_ (.I(_03889_),
    .Z(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08630_ (.I(_03879_),
    .Z(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08631_ (.I0(_03817_),
    .I1(\u2.mem[12][8] ),
    .S(_03890_),
    .Z(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08632_ (.I(_03891_),
    .Z(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08633_ (.I0(_03820_),
    .I1(\u2.mem[12][9] ),
    .S(_03890_),
    .Z(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08634_ (.I(_03892_),
    .Z(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08635_ (.I0(_03822_),
    .I1(\u2.mem[12][10] ),
    .S(_03890_),
    .Z(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08636_ (.I(_03893_),
    .Z(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08637_ (.I0(_03824_),
    .I1(\u2.mem[12][11] ),
    .S(_03890_),
    .Z(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08638_ (.I(_03894_),
    .Z(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08639_ (.I(_03879_),
    .Z(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08640_ (.I0(_03826_),
    .I1(\u2.mem[12][12] ),
    .S(_03895_),
    .Z(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08641_ (.I(_03896_),
    .Z(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08642_ (.I0(_03829_),
    .I1(\u2.mem[12][13] ),
    .S(_03895_),
    .Z(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08643_ (.I(_03897_),
    .Z(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08644_ (.I0(_03831_),
    .I1(\u2.mem[12][14] ),
    .S(_03895_),
    .Z(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08645_ (.I(_03898_),
    .Z(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08646_ (.I0(_03833_),
    .I1(\u2.mem[12][15] ),
    .S(_03895_),
    .Z(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08647_ (.I(_03899_),
    .Z(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08648_ (.I(_03656_),
    .Z(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08649_ (.A1(_03725_),
    .A2(_03482_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08650_ (.A1(_03749_),
    .A2(_03877_),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08651_ (.A1(_03901_),
    .A2(_03902_),
    .ZN(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08652_ (.I(_03903_),
    .Z(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08653_ (.A1(_03480_),
    .A2(_03904_),
    .ZN(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08654_ (.I(_03905_),
    .Z(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08655_ (.I0(_03900_),
    .I1(\u2.mem[13][0] ),
    .S(_03906_),
    .Z(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08656_ (.I(_03907_),
    .Z(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08657_ (.I(_03663_),
    .Z(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08658_ (.I0(_03908_),
    .I1(\u2.mem[13][1] ),
    .S(_03906_),
    .Z(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08659_ (.I(_03909_),
    .Z(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08660_ (.I(_03667_),
    .Z(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08661_ (.I0(_03910_),
    .I1(\u2.mem[13][2] ),
    .S(_03906_),
    .Z(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08662_ (.I(_03911_),
    .Z(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08663_ (.I(_03671_),
    .Z(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08664_ (.I0(_03912_),
    .I1(\u2.mem[13][3] ),
    .S(_03906_),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08665_ (.I(_03913_),
    .Z(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08666_ (.I(_03675_),
    .Z(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08667_ (.I(_03905_),
    .Z(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08668_ (.I0(_03914_),
    .I1(\u2.mem[13][4] ),
    .S(_03915_),
    .Z(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08669_ (.I(_03916_),
    .Z(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08670_ (.I(_03680_),
    .Z(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08671_ (.I0(_03917_),
    .I1(\u2.mem[13][5] ),
    .S(_03915_),
    .Z(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08672_ (.I(_03918_),
    .Z(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08673_ (.I(_03684_),
    .Z(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08674_ (.I0(_03919_),
    .I1(\u2.mem[13][6] ),
    .S(_03915_),
    .Z(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08675_ (.I(_03920_),
    .Z(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08676_ (.I(_03688_),
    .Z(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08677_ (.I0(_03921_),
    .I1(\u2.mem[13][7] ),
    .S(_03915_),
    .Z(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08678_ (.I(_03922_),
    .Z(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08679_ (.I(_03692_),
    .Z(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08680_ (.I(_03905_),
    .Z(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08681_ (.I0(_03923_),
    .I1(\u2.mem[13][8] ),
    .S(_03924_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08682_ (.I(_03925_),
    .Z(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08683_ (.I(_03697_),
    .Z(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08684_ (.I0(_03926_),
    .I1(\u2.mem[13][9] ),
    .S(_03924_),
    .Z(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08685_ (.I(_03927_),
    .Z(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08686_ (.I(_03701_),
    .Z(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08687_ (.I0(_03928_),
    .I1(\u2.mem[13][10] ),
    .S(_03924_),
    .Z(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08688_ (.I(_03929_),
    .Z(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08689_ (.I(_03705_),
    .Z(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08690_ (.I0(_03930_),
    .I1(\u2.mem[13][11] ),
    .S(_03924_),
    .Z(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08691_ (.I(_03931_),
    .Z(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08692_ (.I(_03709_),
    .Z(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08693_ (.I(_03905_),
    .Z(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08694_ (.I0(_03932_),
    .I1(\u2.mem[13][12] ),
    .S(_03933_),
    .Z(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08695_ (.I(_03934_),
    .Z(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08696_ (.I(_03714_),
    .Z(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08697_ (.I0(_03935_),
    .I1(\u2.mem[13][13] ),
    .S(_03933_),
    .Z(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08698_ (.I(_03936_),
    .Z(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08699_ (.I(_03718_),
    .Z(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08700_ (.I0(_03937_),
    .I1(\u2.mem[13][14] ),
    .S(_03933_),
    .Z(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08701_ (.I(_03938_),
    .Z(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08702_ (.I(_03722_),
    .Z(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08703_ (.I0(_03939_),
    .I1(\u2.mem[13][15] ),
    .S(_03933_),
    .Z(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08704_ (.I(_03940_),
    .Z(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08705_ (.A1(_03607_),
    .A2(_03726_),
    .A3(_03878_),
    .ZN(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08706_ (.I(_03941_),
    .Z(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08707_ (.I0(_03900_),
    .I1(\u2.mem[14][0] ),
    .S(_03942_),
    .Z(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08708_ (.I(_03943_),
    .Z(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08709_ (.I0(_03908_),
    .I1(\u2.mem[14][1] ),
    .S(_03942_),
    .Z(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08710_ (.I(_03944_),
    .Z(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08711_ (.I0(_03910_),
    .I1(\u2.mem[14][2] ),
    .S(_03942_),
    .Z(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08712_ (.I(_03945_),
    .Z(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08713_ (.I0(_03912_),
    .I1(\u2.mem[14][3] ),
    .S(_03942_),
    .Z(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08714_ (.I(_03946_),
    .Z(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08715_ (.I(_03941_),
    .Z(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08716_ (.I0(_03914_),
    .I1(\u2.mem[14][4] ),
    .S(_03947_),
    .Z(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08717_ (.I(_03948_),
    .Z(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08718_ (.I0(_03917_),
    .I1(\u2.mem[14][5] ),
    .S(_03947_),
    .Z(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08719_ (.I(_03949_),
    .Z(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08720_ (.I0(_03919_),
    .I1(\u2.mem[14][6] ),
    .S(_03947_),
    .Z(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08721_ (.I(_03950_),
    .Z(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08722_ (.I0(_03921_),
    .I1(\u2.mem[14][7] ),
    .S(_03947_),
    .Z(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08723_ (.I(_03951_),
    .Z(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08724_ (.I(_03941_),
    .Z(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08725_ (.I0(_03923_),
    .I1(\u2.mem[14][8] ),
    .S(_03952_),
    .Z(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08726_ (.I(_03953_),
    .Z(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08727_ (.I0(_03926_),
    .I1(\u2.mem[14][9] ),
    .S(_03952_),
    .Z(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08728_ (.I(_03954_),
    .Z(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08729_ (.I0(_03928_),
    .I1(\u2.mem[14][10] ),
    .S(_03952_),
    .Z(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08730_ (.I(_03955_),
    .Z(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08731_ (.I0(_03930_),
    .I1(\u2.mem[14][11] ),
    .S(_03952_),
    .Z(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08732_ (.I(_03956_),
    .Z(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08733_ (.I(_03941_),
    .Z(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08734_ (.I0(_03932_),
    .I1(\u2.mem[14][12] ),
    .S(_03957_),
    .Z(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08735_ (.I(_03958_),
    .Z(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08736_ (.I0(_03935_),
    .I1(\u2.mem[14][13] ),
    .S(_03957_),
    .Z(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08737_ (.I(_03959_),
    .Z(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08738_ (.I0(_03937_),
    .I1(\u2.mem[14][14] ),
    .S(_03957_),
    .Z(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08739_ (.I(_03960_),
    .Z(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08740_ (.I0(_03939_),
    .I1(\u2.mem[14][15] ),
    .S(_03957_),
    .Z(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08741_ (.I(_03961_),
    .Z(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08742_ (.A1(_03605_),
    .A2(_03606_),
    .A3(_03607_),
    .A4(_03878_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08743_ (.I(_03962_),
    .Z(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08744_ (.I0(_03900_),
    .I1(\u2.mem[15][0] ),
    .S(_03963_),
    .Z(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08745_ (.I(_03964_),
    .Z(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08746_ (.I0(_03908_),
    .I1(\u2.mem[15][1] ),
    .S(_03963_),
    .Z(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08747_ (.I(_03965_),
    .Z(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08748_ (.I0(_03910_),
    .I1(\u2.mem[15][2] ),
    .S(_03963_),
    .Z(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08749_ (.I(_03966_),
    .Z(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08750_ (.I0(_03912_),
    .I1(\u2.mem[15][3] ),
    .S(_03963_),
    .Z(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08751_ (.I(_03967_),
    .Z(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08752_ (.I(_03962_),
    .Z(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08753_ (.I0(_03914_),
    .I1(\u2.mem[15][4] ),
    .S(_03968_),
    .Z(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08754_ (.I(_03969_),
    .Z(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08755_ (.I0(_03917_),
    .I1(\u2.mem[15][5] ),
    .S(_03968_),
    .Z(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08756_ (.I(_03970_),
    .Z(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08757_ (.I0(_03919_),
    .I1(\u2.mem[15][6] ),
    .S(_03968_),
    .Z(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08758_ (.I(_03971_),
    .Z(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08759_ (.I0(_03921_),
    .I1(\u2.mem[15][7] ),
    .S(_03968_),
    .Z(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08760_ (.I(_03972_),
    .Z(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08761_ (.I(_03962_),
    .Z(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08762_ (.I0(_03923_),
    .I1(\u2.mem[15][8] ),
    .S(_03973_),
    .Z(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08763_ (.I(_03974_),
    .Z(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08764_ (.I0(_03926_),
    .I1(\u2.mem[15][9] ),
    .S(_03973_),
    .Z(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08765_ (.I(_03975_),
    .Z(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08766_ (.I0(_03928_),
    .I1(\u2.mem[15][10] ),
    .S(_03973_),
    .Z(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08767_ (.I(_03976_),
    .Z(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08768_ (.I0(_03930_),
    .I1(\u2.mem[15][11] ),
    .S(_03973_),
    .Z(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08769_ (.I(_03977_),
    .Z(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08770_ (.I(_03962_),
    .Z(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08771_ (.I0(_03932_),
    .I1(\u2.mem[15][12] ),
    .S(_03978_),
    .Z(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08772_ (.I(_03979_),
    .Z(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08773_ (.I0(_03935_),
    .I1(\u2.mem[15][13] ),
    .S(_03978_),
    .Z(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08774_ (.I(_03980_),
    .Z(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08775_ (.I0(_03937_),
    .I1(\u2.mem[15][14] ),
    .S(_03978_),
    .Z(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08776_ (.I(_03981_),
    .Z(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08777_ (.I0(_03939_),
    .I1(\u2.mem[15][15] ),
    .S(_03978_),
    .Z(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08778_ (.I(_03982_),
    .Z(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08779_ (.I(_03486_),
    .Z(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08780_ (.I(\mem_address_trans[4].data_sync ),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08781_ (.I(\mem_address_trans[5].data_sync ),
    .Z(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08782_ (.I(\mem_address_trans[7].data_sync ),
    .Z(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08783_ (.A1(_03984_),
    .A2(_03985_),
    .A3(_03478_),
    .A4(_03986_),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08784_ (.I(_03987_),
    .Z(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08785_ (.A1(_03983_),
    .A2(_03988_),
    .ZN(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08786_ (.I(_03989_),
    .Z(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08787_ (.I0(_03900_),
    .I1(\u2.mem[16][0] ),
    .S(_03990_),
    .Z(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08788_ (.I(_03991_),
    .Z(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08789_ (.I0(_03908_),
    .I1(\u2.mem[16][1] ),
    .S(_03990_),
    .Z(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08790_ (.I(_03992_),
    .Z(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08791_ (.I0(_03910_),
    .I1(\u2.mem[16][2] ),
    .S(_03990_),
    .Z(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08792_ (.I(_03993_),
    .Z(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08793_ (.I0(_03912_),
    .I1(\u2.mem[16][3] ),
    .S(_03990_),
    .Z(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08794_ (.I(_03994_),
    .Z(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08795_ (.I(_03989_),
    .Z(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08796_ (.I0(_03914_),
    .I1(\u2.mem[16][4] ),
    .S(_03995_),
    .Z(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08797_ (.I(_03996_),
    .Z(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08798_ (.I0(_03917_),
    .I1(\u2.mem[16][5] ),
    .S(_03995_),
    .Z(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08799_ (.I(_03997_),
    .Z(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08800_ (.I0(_03919_),
    .I1(\u2.mem[16][6] ),
    .S(_03995_),
    .Z(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08801_ (.I(_03998_),
    .Z(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08802_ (.I0(_03921_),
    .I1(\u2.mem[16][7] ),
    .S(_03995_),
    .Z(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08803_ (.I(_03999_),
    .Z(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08804_ (.I(_03989_),
    .Z(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08805_ (.I0(_03923_),
    .I1(\u2.mem[16][8] ),
    .S(_04000_),
    .Z(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08806_ (.I(_04001_),
    .Z(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08807_ (.I0(_03926_),
    .I1(\u2.mem[16][9] ),
    .S(_04000_),
    .Z(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08808_ (.I(_04002_),
    .Z(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08809_ (.I0(_03928_),
    .I1(\u2.mem[16][10] ),
    .S(_04000_),
    .Z(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08810_ (.I(_04003_),
    .Z(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08811_ (.I0(_03930_),
    .I1(\u2.mem[16][11] ),
    .S(_04000_),
    .Z(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08812_ (.I(_04004_),
    .Z(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08813_ (.I(_03989_),
    .Z(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08814_ (.I0(_03932_),
    .I1(\u2.mem[16][12] ),
    .S(_04005_),
    .Z(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08815_ (.I(_04006_),
    .Z(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08816_ (.I0(_03935_),
    .I1(\u2.mem[16][13] ),
    .S(_04005_),
    .Z(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08817_ (.I(_04007_),
    .Z(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08818_ (.I0(_03937_),
    .I1(\u2.mem[16][14] ),
    .S(_04005_),
    .Z(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08819_ (.I(_04008_),
    .Z(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08820_ (.I0(_03939_),
    .I1(\u2.mem[16][15] ),
    .S(_04005_),
    .Z(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08821_ (.I(_04009_),
    .Z(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08822_ (.I(_03656_),
    .Z(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08823_ (.I(_03987_),
    .Z(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08824_ (.A1(_03483_),
    .A2(_03540_),
    .A3(_03544_),
    .Z(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08825_ (.I(_04012_),
    .Z(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08826_ (.A1(_04011_),
    .A2(_04013_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08827_ (.I(_04014_),
    .Z(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08828_ (.I0(_04010_),
    .I1(\u2.mem[17][0] ),
    .S(_04015_),
    .Z(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08829_ (.I(_04016_),
    .Z(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08830_ (.I(_03663_),
    .Z(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08831_ (.I0(_04017_),
    .I1(\u2.mem[17][1] ),
    .S(_04015_),
    .Z(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08832_ (.I(_04018_),
    .Z(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08833_ (.I(_03667_),
    .Z(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08834_ (.I0(_04019_),
    .I1(\u2.mem[17][2] ),
    .S(_04015_),
    .Z(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08835_ (.I(_04020_),
    .Z(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08836_ (.I(_03671_),
    .Z(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08837_ (.I0(_04021_),
    .I1(\u2.mem[17][3] ),
    .S(_04015_),
    .Z(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08838_ (.I(_04022_),
    .Z(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08839_ (.I(_03675_),
    .Z(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08840_ (.I(_04014_),
    .Z(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08841_ (.I0(_04023_),
    .I1(\u2.mem[17][4] ),
    .S(_04024_),
    .Z(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08842_ (.I(_04025_),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08843_ (.I(_03680_),
    .Z(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08844_ (.I0(_04026_),
    .I1(\u2.mem[17][5] ),
    .S(_04024_),
    .Z(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08845_ (.I(_04027_),
    .Z(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08846_ (.I(_03684_),
    .Z(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08847_ (.I0(_04028_),
    .I1(\u2.mem[17][6] ),
    .S(_04024_),
    .Z(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08848_ (.I(_04029_),
    .Z(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08849_ (.I(_03688_),
    .Z(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08850_ (.I0(_04030_),
    .I1(\u2.mem[17][7] ),
    .S(_04024_),
    .Z(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08851_ (.I(_04031_),
    .Z(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08852_ (.I(_03692_),
    .Z(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08853_ (.I(_04014_),
    .Z(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08854_ (.I0(_04032_),
    .I1(\u2.mem[17][8] ),
    .S(_04033_),
    .Z(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08855_ (.I(_04034_),
    .Z(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08856_ (.I(_03697_),
    .Z(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08857_ (.I0(_04035_),
    .I1(\u2.mem[17][9] ),
    .S(_04033_),
    .Z(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08858_ (.I(_04036_),
    .Z(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08859_ (.I(_03701_),
    .Z(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08860_ (.I0(_04037_),
    .I1(\u2.mem[17][10] ),
    .S(_04033_),
    .Z(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08861_ (.I(_04038_),
    .Z(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08862_ (.I(_03705_),
    .Z(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08863_ (.I0(_04039_),
    .I1(\u2.mem[17][11] ),
    .S(_04033_),
    .Z(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08864_ (.I(_04040_),
    .Z(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08865_ (.I(_03709_),
    .Z(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08866_ (.I(_04014_),
    .Z(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08867_ (.I0(_04041_),
    .I1(\u2.mem[17][12] ),
    .S(_04042_),
    .Z(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08868_ (.I(_04043_),
    .Z(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08869_ (.I(_03714_),
    .Z(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08870_ (.I0(_04044_),
    .I1(\u2.mem[17][13] ),
    .S(_04042_),
    .Z(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08871_ (.I(_04045_),
    .Z(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08872_ (.I(_03718_),
    .Z(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08873_ (.I0(_04046_),
    .I1(\u2.mem[17][14] ),
    .S(_04042_),
    .Z(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08874_ (.I(_04047_),
    .Z(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08875_ (.I(_03722_),
    .Z(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08876_ (.I0(_04048_),
    .I1(\u2.mem[17][15] ),
    .S(_04042_),
    .Z(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08877_ (.I(_04049_),
    .Z(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08878_ (.A1(_03583_),
    .A2(_03988_),
    .ZN(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08879_ (.I(_04050_),
    .Z(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08880_ (.I0(_04010_),
    .I1(\u2.mem[18][0] ),
    .S(_04051_),
    .Z(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08881_ (.I(_04052_),
    .Z(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08882_ (.I0(_04017_),
    .I1(\u2.mem[18][1] ),
    .S(_04051_),
    .Z(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08883_ (.I(_04053_),
    .Z(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08884_ (.I0(_04019_),
    .I1(\u2.mem[18][2] ),
    .S(_04051_),
    .Z(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08885_ (.I(_04054_),
    .Z(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08886_ (.I0(_04021_),
    .I1(\u2.mem[18][3] ),
    .S(_04051_),
    .Z(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08887_ (.I(_04055_),
    .Z(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08888_ (.I(_04050_),
    .Z(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08889_ (.I0(_04023_),
    .I1(\u2.mem[18][4] ),
    .S(_04056_),
    .Z(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08890_ (.I(_04057_),
    .Z(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08891_ (.I0(_04026_),
    .I1(\u2.mem[18][5] ),
    .S(_04056_),
    .Z(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08892_ (.I(_04058_),
    .Z(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08893_ (.I0(_04028_),
    .I1(\u2.mem[18][6] ),
    .S(_04056_),
    .Z(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08894_ (.I(_04059_),
    .Z(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08895_ (.I0(_04030_),
    .I1(\u2.mem[18][7] ),
    .S(_04056_),
    .Z(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08896_ (.I(_04060_),
    .Z(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08897_ (.I(_04050_),
    .Z(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08898_ (.I0(_04032_),
    .I1(\u2.mem[18][8] ),
    .S(_04061_),
    .Z(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08899_ (.I(_04062_),
    .Z(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08900_ (.I0(_04035_),
    .I1(\u2.mem[18][9] ),
    .S(_04061_),
    .Z(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08901_ (.I(_04063_),
    .Z(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08902_ (.I0(_04037_),
    .I1(\u2.mem[18][10] ),
    .S(_04061_),
    .Z(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08903_ (.I(_04064_),
    .Z(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08904_ (.I0(_04039_),
    .I1(\u2.mem[18][11] ),
    .S(_04061_),
    .Z(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08905_ (.I(_04065_),
    .Z(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08906_ (.I(_04050_),
    .Z(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08907_ (.I0(_04041_),
    .I1(\u2.mem[18][12] ),
    .S(_04066_),
    .Z(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08908_ (.I(_04067_),
    .Z(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08909_ (.I0(_04044_),
    .I1(\u2.mem[18][13] ),
    .S(_04066_),
    .Z(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08910_ (.I(_04068_),
    .Z(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08911_ (.I0(_04046_),
    .I1(\u2.mem[18][14] ),
    .S(_04066_),
    .Z(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08912_ (.I(_04069_),
    .Z(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08913_ (.I0(_04048_),
    .I1(\u2.mem[18][15] ),
    .S(_04066_),
    .Z(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08914_ (.I(_04070_),
    .Z(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08915_ (.A1(_03485_),
    .A2(_03748_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08916_ (.I(_04071_),
    .Z(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08917_ (.A1(_04072_),
    .A2(_03988_),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08918_ (.I(_04073_),
    .Z(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08919_ (.I0(_04010_),
    .I1(\u2.mem[19][0] ),
    .S(_04074_),
    .Z(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08920_ (.I(_04075_),
    .Z(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08921_ (.I0(_04017_),
    .I1(\u2.mem[19][1] ),
    .S(_04074_),
    .Z(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08922_ (.I(_04076_),
    .Z(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08923_ (.I0(_04019_),
    .I1(\u2.mem[19][2] ),
    .S(_04074_),
    .Z(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08924_ (.I(_04077_),
    .Z(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08925_ (.I0(_04021_),
    .I1(\u2.mem[19][3] ),
    .S(_04074_),
    .Z(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08926_ (.I(_04078_),
    .Z(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08927_ (.I(_04073_),
    .Z(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08928_ (.I0(_04023_),
    .I1(\u2.mem[19][4] ),
    .S(_04079_),
    .Z(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08929_ (.I(_04080_),
    .Z(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08930_ (.I0(_04026_),
    .I1(\u2.mem[19][5] ),
    .S(_04079_),
    .Z(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08931_ (.I(_04081_),
    .Z(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08932_ (.I0(_04028_),
    .I1(\u2.mem[19][6] ),
    .S(_04079_),
    .Z(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08933_ (.I(_04082_),
    .Z(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08934_ (.I0(_04030_),
    .I1(\u2.mem[19][7] ),
    .S(_04079_),
    .Z(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08935_ (.I(_04083_),
    .Z(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08936_ (.I(_04073_),
    .Z(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08937_ (.I0(_04032_),
    .I1(\u2.mem[19][8] ),
    .S(_04084_),
    .Z(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08938_ (.I(_04085_),
    .Z(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08939_ (.I0(_04035_),
    .I1(\u2.mem[19][9] ),
    .S(_04084_),
    .Z(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08940_ (.I(_04086_),
    .Z(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08941_ (.I0(_04037_),
    .I1(\u2.mem[19][10] ),
    .S(_04084_),
    .Z(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08942_ (.I(_04087_),
    .Z(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08943_ (.I0(_04039_),
    .I1(\u2.mem[19][11] ),
    .S(_04084_),
    .Z(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08944_ (.I(_04088_),
    .Z(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08945_ (.I(_04073_),
    .Z(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08946_ (.I0(_04041_),
    .I1(\u2.mem[19][12] ),
    .S(_04089_),
    .Z(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08947_ (.I(_04090_),
    .Z(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08948_ (.I0(_04044_),
    .I1(\u2.mem[19][13] ),
    .S(_04089_),
    .Z(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08949_ (.I(_04091_),
    .Z(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08950_ (.I0(_04046_),
    .I1(\u2.mem[19][14] ),
    .S(_04089_),
    .Z(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08951_ (.I(_04092_),
    .Z(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08952_ (.I0(_04048_),
    .I1(\u2.mem[19][15] ),
    .S(_04089_),
    .Z(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08953_ (.I(_04093_),
    .Z(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _08954_ (.A1(_03629_),
    .A2(_03540_),
    .A3(_03633_),
    .Z(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08955_ (.I(_04094_),
    .Z(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08956_ (.A1(_04095_),
    .A2(_03988_),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08957_ (.I(_04096_),
    .Z(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08958_ (.I0(_04010_),
    .I1(\u2.mem[20][0] ),
    .S(_04097_),
    .Z(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08959_ (.I(_04098_),
    .Z(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08960_ (.I0(_04017_),
    .I1(\u2.mem[20][1] ),
    .S(_04097_),
    .Z(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08961_ (.I(_04099_),
    .Z(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08962_ (.I0(_04019_),
    .I1(\u2.mem[20][2] ),
    .S(_04097_),
    .Z(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08963_ (.I(_04100_),
    .Z(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08964_ (.I0(_04021_),
    .I1(\u2.mem[20][3] ),
    .S(_04097_),
    .Z(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08965_ (.I(_04101_),
    .Z(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08966_ (.I(_04096_),
    .Z(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08967_ (.I0(_04023_),
    .I1(\u2.mem[20][4] ),
    .S(_04102_),
    .Z(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08968_ (.I(_04103_),
    .Z(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08969_ (.I0(_04026_),
    .I1(\u2.mem[20][5] ),
    .S(_04102_),
    .Z(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08970_ (.I(_04104_),
    .Z(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08971_ (.I0(_04028_),
    .I1(\u2.mem[20][6] ),
    .S(_04102_),
    .Z(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08972_ (.I(_04105_),
    .Z(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08973_ (.I0(_04030_),
    .I1(\u2.mem[20][7] ),
    .S(_04102_),
    .Z(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08974_ (.I(_04106_),
    .Z(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08975_ (.I(_04096_),
    .Z(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08976_ (.I0(_04032_),
    .I1(\u2.mem[20][8] ),
    .S(_04107_),
    .Z(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08977_ (.I(_04108_),
    .Z(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08978_ (.I0(_04035_),
    .I1(\u2.mem[20][9] ),
    .S(_04107_),
    .Z(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08979_ (.I(_04109_),
    .Z(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08980_ (.I0(_04037_),
    .I1(\u2.mem[20][10] ),
    .S(_04107_),
    .Z(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08981_ (.I(_04110_),
    .Z(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08982_ (.I0(_04039_),
    .I1(\u2.mem[20][11] ),
    .S(_04107_),
    .Z(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08983_ (.I(_04111_),
    .Z(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08984_ (.I(_04096_),
    .Z(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08985_ (.I0(_04041_),
    .I1(\u2.mem[20][12] ),
    .S(_04112_),
    .Z(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08986_ (.I(_04113_),
    .Z(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08987_ (.I0(_04044_),
    .I1(\u2.mem[20][13] ),
    .S(_04112_),
    .Z(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08988_ (.I(_04114_),
    .Z(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08989_ (.I0(_04046_),
    .I1(\u2.mem[20][14] ),
    .S(_04112_),
    .Z(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08990_ (.I(_04115_),
    .Z(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08991_ (.I0(_04048_),
    .I1(\u2.mem[20][15] ),
    .S(_04112_),
    .Z(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08992_ (.I(_04116_),
    .Z(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08993_ (.I(\data_in_trans[0].data_sync ),
    .Z(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08994_ (.I(_04117_),
    .Z(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08995_ (.I(_04118_),
    .Z(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08996_ (.A1(_03901_),
    .A2(_03750_),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08997_ (.I(_04120_),
    .Z(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08998_ (.I(_03987_),
    .Z(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08999_ (.A1(_04121_),
    .A2(_04122_),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09000_ (.I(_04123_),
    .Z(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09001_ (.I0(_04119_),
    .I1(\u2.mem[21][0] ),
    .S(_04124_),
    .Z(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09002_ (.I(_04125_),
    .Z(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09003_ (.I(\data_in_trans[1].data_sync ),
    .Z(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09004_ (.I(_04126_),
    .Z(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09005_ (.I(_04127_),
    .Z(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09006_ (.I0(_04128_),
    .I1(\u2.mem[21][1] ),
    .S(_04124_),
    .Z(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09007_ (.I(_04129_),
    .Z(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09008_ (.I(\data_in_trans[2].data_sync ),
    .Z(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09009_ (.I(_04130_),
    .Z(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09010_ (.I(_04131_),
    .Z(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09011_ (.I0(_04132_),
    .I1(\u2.mem[21][2] ),
    .S(_04124_),
    .Z(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09012_ (.I(_04133_),
    .Z(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09013_ (.I(\data_in_trans[3].data_sync ),
    .Z(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09014_ (.I(_04134_),
    .Z(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09015_ (.I(_04135_),
    .Z(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09016_ (.I0(_04136_),
    .I1(\u2.mem[21][3] ),
    .S(_04124_),
    .Z(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09017_ (.I(_04137_),
    .Z(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09018_ (.I(\data_in_trans[4].data_sync ),
    .Z(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09019_ (.I(_04138_),
    .Z(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09020_ (.I(_04139_),
    .Z(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09021_ (.I(_04123_),
    .Z(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09022_ (.I0(_04140_),
    .I1(\u2.mem[21][4] ),
    .S(_04141_),
    .Z(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09023_ (.I(_04142_),
    .Z(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09024_ (.I(\data_in_trans[5].data_sync ),
    .Z(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09025_ (.I(_04143_),
    .Z(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09026_ (.I(_04144_),
    .Z(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09027_ (.I0(_04145_),
    .I1(\u2.mem[21][5] ),
    .S(_04141_),
    .Z(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09028_ (.I(_04146_),
    .Z(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09029_ (.I(\data_in_trans[6].data_sync ),
    .Z(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09030_ (.I(_04147_),
    .Z(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09031_ (.I0(_04148_),
    .I1(\u2.mem[21][6] ),
    .S(_04141_),
    .Z(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09032_ (.I(_04149_),
    .Z(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09033_ (.I(\data_in_trans[7].data_sync ),
    .Z(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09034_ (.I(_04150_),
    .Z(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09035_ (.I0(_04151_),
    .I1(\u2.mem[21][7] ),
    .S(_04141_),
    .Z(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09036_ (.I(_04152_),
    .Z(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09037_ (.I(\data_in_trans[8].data_sync ),
    .Z(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09038_ (.I(_04153_),
    .Z(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09039_ (.I(_04123_),
    .Z(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09040_ (.I0(_04154_),
    .I1(\u2.mem[21][8] ),
    .S(_04155_),
    .Z(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09041_ (.I(_04156_),
    .Z(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09042_ (.I(\data_in_trans[9].data_sync ),
    .Z(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09043_ (.I(_04157_),
    .Z(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09044_ (.I0(_04158_),
    .I1(\u2.mem[21][9] ),
    .S(_04155_),
    .Z(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09045_ (.I(_04159_),
    .Z(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09046_ (.I(\data_in_trans[10].data_sync ),
    .Z(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09047_ (.I(_04160_),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09048_ (.I0(_04161_),
    .I1(\u2.mem[21][10] ),
    .S(_04155_),
    .Z(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09049_ (.I(_04162_),
    .Z(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09050_ (.I(\data_in_trans[11].data_sync ),
    .Z(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09051_ (.I(_04163_),
    .Z(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09052_ (.I0(_04164_),
    .I1(\u2.mem[21][11] ),
    .S(_04155_),
    .Z(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09053_ (.I(_04165_),
    .Z(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09054_ (.I(\data_in_trans[12].data_sync ),
    .Z(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09055_ (.I(_04166_),
    .Z(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09056_ (.I(_04123_),
    .Z(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09057_ (.I0(_04167_),
    .I1(\u2.mem[21][12] ),
    .S(_04168_),
    .Z(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09058_ (.I(_04169_),
    .Z(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09059_ (.I(\data_in_trans[13].data_sync ),
    .Z(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09060_ (.I(_04170_),
    .Z(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09061_ (.I0(_04171_),
    .I1(\u2.mem[21][13] ),
    .S(_04168_),
    .Z(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09062_ (.I(_04172_),
    .Z(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09063_ (.I(\data_in_trans[14].data_sync ),
    .Z(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09064_ (.I(_04173_),
    .Z(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09065_ (.I0(_04174_),
    .I1(\u2.mem[21][14] ),
    .S(_04168_),
    .Z(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09066_ (.I(_04175_),
    .Z(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09067_ (.I(\data_in_trans[15].data_sync ),
    .Z(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09068_ (.I(_04176_),
    .Z(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09069_ (.I0(_04177_),
    .I1(\u2.mem[21][15] ),
    .S(_04168_),
    .Z(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09070_ (.I(_04178_),
    .Z(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09071_ (.A1(_03581_),
    .A2(_03750_),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09072_ (.I(_04179_),
    .Z(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09073_ (.A1(_04180_),
    .A2(_04122_),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09074_ (.I(_04181_),
    .Z(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09075_ (.I0(_04119_),
    .I1(\u2.mem[22][0] ),
    .S(_04182_),
    .Z(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09076_ (.I(_04183_),
    .Z(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09077_ (.I0(_04128_),
    .I1(\u2.mem[22][1] ),
    .S(_04182_),
    .Z(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09078_ (.I(_04184_),
    .Z(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09079_ (.I0(_04132_),
    .I1(\u2.mem[22][2] ),
    .S(_04182_),
    .Z(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09080_ (.I(_04185_),
    .Z(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09081_ (.I0(_04136_),
    .I1(\u2.mem[22][3] ),
    .S(_04182_),
    .Z(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09082_ (.I(_04186_),
    .Z(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09083_ (.I(_04181_),
    .Z(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09084_ (.I0(_04140_),
    .I1(\u2.mem[22][4] ),
    .S(_04187_),
    .Z(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09085_ (.I(_04188_),
    .Z(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09086_ (.I0(_04145_),
    .I1(\u2.mem[22][5] ),
    .S(_04187_),
    .Z(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09087_ (.I(_04189_),
    .Z(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09088_ (.I0(_04148_),
    .I1(\u2.mem[22][6] ),
    .S(_04187_),
    .Z(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09089_ (.I(_04190_),
    .Z(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09090_ (.I0(_04151_),
    .I1(\u2.mem[22][7] ),
    .S(_04187_),
    .Z(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09091_ (.I(_04191_),
    .Z(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09092_ (.I(_04181_),
    .Z(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09093_ (.I0(_04154_),
    .I1(\u2.mem[22][8] ),
    .S(_04192_),
    .Z(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09094_ (.I(_04193_),
    .Z(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09095_ (.I0(_04158_),
    .I1(\u2.mem[22][9] ),
    .S(_04192_),
    .Z(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09096_ (.I(_04194_),
    .Z(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09097_ (.I0(_04161_),
    .I1(\u2.mem[22][10] ),
    .S(_04192_),
    .Z(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09098_ (.I(_04195_),
    .Z(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09099_ (.I0(_04164_),
    .I1(\u2.mem[22][11] ),
    .S(_04192_),
    .Z(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09100_ (.I(_04196_),
    .Z(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09101_ (.I(_04181_),
    .Z(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09102_ (.I0(_04167_),
    .I1(\u2.mem[22][12] ),
    .S(_04197_),
    .Z(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09103_ (.I(_04198_),
    .Z(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09104_ (.I0(_04171_),
    .I1(\u2.mem[22][13] ),
    .S(_04197_),
    .Z(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09105_ (.I(_04199_),
    .Z(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09106_ (.I0(_04174_),
    .I1(\u2.mem[22][14] ),
    .S(_04197_),
    .Z(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09107_ (.I(_04200_),
    .Z(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09108_ (.I0(_04177_),
    .I1(\u2.mem[22][15] ),
    .S(_04197_),
    .Z(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09109_ (.I(_04201_),
    .Z(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09110_ (.A1(_03752_),
    .A2(_04122_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09111_ (.I(_04202_),
    .Z(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09112_ (.I0(_04119_),
    .I1(\u2.mem[23][0] ),
    .S(_04203_),
    .Z(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09113_ (.I(_04204_),
    .Z(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09114_ (.I0(_04128_),
    .I1(\u2.mem[23][1] ),
    .S(_04203_),
    .Z(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09115_ (.I(_04205_),
    .Z(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09116_ (.I0(_04132_),
    .I1(\u2.mem[23][2] ),
    .S(_04203_),
    .Z(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09117_ (.I(_04206_),
    .Z(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09118_ (.I0(_04136_),
    .I1(\u2.mem[23][3] ),
    .S(_04203_),
    .Z(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09119_ (.I(_04207_),
    .Z(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09120_ (.I(_04202_),
    .Z(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09121_ (.I0(_04140_),
    .I1(\u2.mem[23][4] ),
    .S(_04208_),
    .Z(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09122_ (.I(_04209_),
    .Z(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09123_ (.I0(_04145_),
    .I1(\u2.mem[23][5] ),
    .S(_04208_),
    .Z(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09124_ (.I(_04210_),
    .Z(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09125_ (.I0(_04148_),
    .I1(\u2.mem[23][6] ),
    .S(_04208_),
    .Z(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09126_ (.I(_04211_),
    .Z(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09127_ (.I0(_04151_),
    .I1(\u2.mem[23][7] ),
    .S(_04208_),
    .Z(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09128_ (.I(_04212_),
    .Z(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09129_ (.I(_04202_),
    .Z(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09130_ (.I0(_04154_),
    .I1(\u2.mem[23][8] ),
    .S(_04213_),
    .Z(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09131_ (.I(_04214_),
    .Z(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09132_ (.I0(_04158_),
    .I1(\u2.mem[23][9] ),
    .S(_04213_),
    .Z(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09133_ (.I(_04215_),
    .Z(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09134_ (.I0(_04161_),
    .I1(\u2.mem[23][10] ),
    .S(_04213_),
    .Z(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09135_ (.I(_04216_),
    .Z(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09136_ (.I0(_04164_),
    .I1(\u2.mem[23][11] ),
    .S(_04213_),
    .Z(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09137_ (.I(_04217_),
    .Z(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09138_ (.I(_04202_),
    .Z(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09139_ (.I0(_04167_),
    .I1(\u2.mem[23][12] ),
    .S(_04218_),
    .Z(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09140_ (.I(_04219_),
    .Z(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09141_ (.I0(_04171_),
    .I1(\u2.mem[23][13] ),
    .S(_04218_),
    .Z(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09142_ (.I(_04220_),
    .Z(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09143_ (.I0(_04174_),
    .I1(\u2.mem[23][14] ),
    .S(_04218_),
    .Z(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09144_ (.I(_04221_),
    .Z(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09145_ (.I0(_04177_),
    .I1(\u2.mem[23][15] ),
    .S(_04218_),
    .Z(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09146_ (.I(_04222_),
    .Z(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _09147_ (.A1(_03629_),
    .A2(_03749_),
    .A3(_03775_),
    .Z(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09148_ (.I(_04223_),
    .Z(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09149_ (.A1(_04224_),
    .A2(_04122_),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09150_ (.I(_04225_),
    .Z(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09151_ (.I0(_04119_),
    .I1(\u2.mem[24][0] ),
    .S(_04226_),
    .Z(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09152_ (.I(_04227_),
    .Z(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09153_ (.I0(_04128_),
    .I1(\u2.mem[24][1] ),
    .S(_04226_),
    .Z(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09154_ (.I(_04228_),
    .Z(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09155_ (.I0(_04132_),
    .I1(\u2.mem[24][2] ),
    .S(_04226_),
    .Z(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09156_ (.I(_04229_),
    .Z(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09157_ (.I0(_04136_),
    .I1(\u2.mem[24][3] ),
    .S(_04226_),
    .Z(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09158_ (.I(_04230_),
    .Z(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09159_ (.I(_04225_),
    .Z(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09160_ (.I0(_04140_),
    .I1(\u2.mem[24][4] ),
    .S(_04231_),
    .Z(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09161_ (.I(_04232_),
    .Z(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09162_ (.I0(_04145_),
    .I1(\u2.mem[24][5] ),
    .S(_04231_),
    .Z(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09163_ (.I(_04233_),
    .Z(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09164_ (.I0(_04148_),
    .I1(\u2.mem[24][6] ),
    .S(_04231_),
    .Z(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09165_ (.I(_04234_),
    .Z(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09166_ (.I0(_04151_),
    .I1(\u2.mem[24][7] ),
    .S(_04231_),
    .Z(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09167_ (.I(_04235_),
    .Z(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09168_ (.I(_04225_),
    .Z(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09169_ (.I0(_04154_),
    .I1(\u2.mem[24][8] ),
    .S(_04236_),
    .Z(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09170_ (.I(_04237_),
    .Z(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09171_ (.I0(_04158_),
    .I1(\u2.mem[24][9] ),
    .S(_04236_),
    .Z(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09172_ (.I(_04238_),
    .Z(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09173_ (.I0(_04161_),
    .I1(\u2.mem[24][10] ),
    .S(_04236_),
    .Z(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09174_ (.I(_04239_),
    .Z(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09175_ (.I0(_04164_),
    .I1(\u2.mem[24][11] ),
    .S(_04236_),
    .Z(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09176_ (.I(_04240_),
    .Z(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09177_ (.I(_04225_),
    .Z(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09178_ (.I0(_04167_),
    .I1(\u2.mem[24][12] ),
    .S(_04241_),
    .Z(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09179_ (.I(_04242_),
    .Z(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09180_ (.I0(_04171_),
    .I1(\u2.mem[24][13] ),
    .S(_04241_),
    .Z(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09181_ (.I(_04243_),
    .Z(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09182_ (.I0(_04174_),
    .I1(\u2.mem[24][14] ),
    .S(_04241_),
    .Z(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09183_ (.I(_04244_),
    .Z(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09184_ (.I0(_04177_),
    .I1(\u2.mem[24][15] ),
    .S(_04241_),
    .Z(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09185_ (.I(_04245_),
    .Z(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09186_ (.I(_04118_),
    .Z(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09187_ (.A1(_03749_),
    .A2(_03775_),
    .ZN(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09188_ (.A1(_03901_),
    .A2(_04247_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09189_ (.I(_04248_),
    .Z(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09190_ (.I(_03987_),
    .Z(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09191_ (.A1(_04249_),
    .A2(_04250_),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09192_ (.I(_04251_),
    .Z(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09193_ (.I0(_04246_),
    .I1(\u2.mem[25][0] ),
    .S(_04252_),
    .Z(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09194_ (.I(_04253_),
    .Z(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09195_ (.I(_04127_),
    .Z(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09196_ (.I0(_04254_),
    .I1(\u2.mem[25][1] ),
    .S(_04252_),
    .Z(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09197_ (.I(_04255_),
    .Z(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09198_ (.I(_04131_),
    .Z(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09199_ (.I0(_04256_),
    .I1(\u2.mem[25][2] ),
    .S(_04252_),
    .Z(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09200_ (.I(_04257_),
    .Z(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09201_ (.I(_04135_),
    .Z(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09202_ (.I0(_04258_),
    .I1(\u2.mem[25][3] ),
    .S(_04252_),
    .Z(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09203_ (.I(_04259_),
    .Z(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09204_ (.I(_04139_),
    .Z(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09205_ (.I(_04251_),
    .Z(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09206_ (.I0(_04260_),
    .I1(\u2.mem[25][4] ),
    .S(_04261_),
    .Z(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09207_ (.I(_04262_),
    .Z(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09208_ (.I(_04144_),
    .Z(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09209_ (.I0(_04263_),
    .I1(\u2.mem[25][5] ),
    .S(_04261_),
    .Z(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09210_ (.I(_04264_),
    .Z(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09211_ (.I(_04147_),
    .Z(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09212_ (.I0(_04265_),
    .I1(\u2.mem[25][6] ),
    .S(_04261_),
    .Z(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09213_ (.I(_04266_),
    .Z(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09214_ (.I(_04150_),
    .Z(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09215_ (.I0(_04267_),
    .I1(\u2.mem[25][7] ),
    .S(_04261_),
    .Z(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09216_ (.I(_04268_),
    .Z(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09217_ (.I(_04153_),
    .Z(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09218_ (.I(_04251_),
    .Z(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09219_ (.I0(_04269_),
    .I1(\u2.mem[25][8] ),
    .S(_04270_),
    .Z(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09220_ (.I(_04271_),
    .Z(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09221_ (.I(_04157_),
    .Z(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09222_ (.I0(_04272_),
    .I1(\u2.mem[25][9] ),
    .S(_04270_),
    .Z(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09223_ (.I(_04273_),
    .Z(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09224_ (.I(_04160_),
    .Z(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09225_ (.I0(_04274_),
    .I1(\u2.mem[25][10] ),
    .S(_04270_),
    .Z(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09226_ (.I(_04275_),
    .Z(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09227_ (.I(_04163_),
    .Z(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09228_ (.I0(_04276_),
    .I1(\u2.mem[25][11] ),
    .S(_04270_),
    .Z(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09229_ (.I(_04277_),
    .Z(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09230_ (.I(_04166_),
    .Z(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09231_ (.I(_04251_),
    .Z(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09232_ (.I0(_04278_),
    .I1(\u2.mem[25][12] ),
    .S(_04279_),
    .Z(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09233_ (.I(_04280_),
    .Z(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09234_ (.I(_04170_),
    .Z(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09235_ (.I0(_04281_),
    .I1(\u2.mem[25][13] ),
    .S(_04279_),
    .Z(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09236_ (.I(_04282_),
    .Z(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09237_ (.I(_04173_),
    .Z(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09238_ (.I0(_04283_),
    .I1(\u2.mem[25][14] ),
    .S(_04279_),
    .Z(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09239_ (.I(_04284_),
    .Z(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09240_ (.I(_04176_),
    .Z(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09241_ (.I0(_04285_),
    .I1(\u2.mem[25][15] ),
    .S(_04279_),
    .Z(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09242_ (.I(_04286_),
    .Z(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09243_ (.A1(_03581_),
    .A2(_04247_),
    .ZN(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09244_ (.I(_04287_),
    .Z(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09245_ (.A1(_04288_),
    .A2(_04250_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09246_ (.I(_04289_),
    .Z(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09247_ (.I0(_04246_),
    .I1(\u2.mem[26][0] ),
    .S(_04290_),
    .Z(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09248_ (.I(_04291_),
    .Z(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09249_ (.I0(_04254_),
    .I1(\u2.mem[26][1] ),
    .S(_04290_),
    .Z(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09250_ (.I(_04292_),
    .Z(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09251_ (.I0(_04256_),
    .I1(\u2.mem[26][2] ),
    .S(_04290_),
    .Z(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09252_ (.I(_04293_),
    .Z(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09253_ (.I0(_04258_),
    .I1(\u2.mem[26][3] ),
    .S(_04290_),
    .Z(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09254_ (.I(_04294_),
    .Z(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09255_ (.I(_04289_),
    .Z(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09256_ (.I0(_04260_),
    .I1(\u2.mem[26][4] ),
    .S(_04295_),
    .Z(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09257_ (.I(_04296_),
    .Z(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09258_ (.I0(_04263_),
    .I1(\u2.mem[26][5] ),
    .S(_04295_),
    .Z(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09259_ (.I(_04297_),
    .Z(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09260_ (.I0(_04265_),
    .I1(\u2.mem[26][6] ),
    .S(_04295_),
    .Z(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09261_ (.I(_04298_),
    .Z(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09262_ (.I0(_04267_),
    .I1(\u2.mem[26][7] ),
    .S(_04295_),
    .Z(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09263_ (.I(_04299_),
    .Z(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09264_ (.I(_04289_),
    .Z(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09265_ (.I0(_04269_),
    .I1(\u2.mem[26][8] ),
    .S(_04300_),
    .Z(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09266_ (.I(_04301_),
    .Z(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09267_ (.I0(_04272_),
    .I1(\u2.mem[26][9] ),
    .S(_04300_),
    .Z(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09268_ (.I(_04302_),
    .Z(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09269_ (.I0(_04274_),
    .I1(\u2.mem[26][10] ),
    .S(_04300_),
    .Z(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09270_ (.I(_04303_),
    .Z(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09271_ (.I0(_04276_),
    .I1(\u2.mem[26][11] ),
    .S(_04300_),
    .Z(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09272_ (.I(_04304_),
    .Z(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09273_ (.I(_04289_),
    .Z(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09274_ (.I0(_04278_),
    .I1(\u2.mem[26][12] ),
    .S(_04305_),
    .Z(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09275_ (.I(_04306_),
    .Z(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09276_ (.I0(_04281_),
    .I1(\u2.mem[26][13] ),
    .S(_04305_),
    .Z(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09277_ (.I(_04307_),
    .Z(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09278_ (.I0(_04283_),
    .I1(\u2.mem[26][14] ),
    .S(_04305_),
    .Z(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09279_ (.I(_04308_),
    .Z(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09280_ (.I0(_04285_),
    .I1(\u2.mem[26][15] ),
    .S(_04305_),
    .Z(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09281_ (.I(_04309_),
    .Z(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09282_ (.A1(_03748_),
    .A2(_04247_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09283_ (.I(_04310_),
    .Z(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09284_ (.A1(_04311_),
    .A2(_04250_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09285_ (.I(_04312_),
    .Z(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09286_ (.I0(_04246_),
    .I1(\u2.mem[27][0] ),
    .S(_04313_),
    .Z(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09287_ (.I(_04314_),
    .Z(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09288_ (.I0(_04254_),
    .I1(\u2.mem[27][1] ),
    .S(_04313_),
    .Z(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09289_ (.I(_04315_),
    .Z(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09290_ (.I0(_04256_),
    .I1(\u2.mem[27][2] ),
    .S(_04313_),
    .Z(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09291_ (.I(_04316_),
    .Z(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09292_ (.I0(_04258_),
    .I1(\u2.mem[27][3] ),
    .S(_04313_),
    .Z(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09293_ (.I(_04317_),
    .Z(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09294_ (.I(_04312_),
    .Z(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09295_ (.I0(_04260_),
    .I1(\u2.mem[27][4] ),
    .S(_04318_),
    .Z(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09296_ (.I(_04319_),
    .Z(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09297_ (.I0(_04263_),
    .I1(\u2.mem[27][5] ),
    .S(_04318_),
    .Z(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09298_ (.I(_04320_),
    .Z(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09299_ (.I0(_04265_),
    .I1(\u2.mem[27][6] ),
    .S(_04318_),
    .Z(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09300_ (.I(_04321_),
    .Z(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09301_ (.I0(_04267_),
    .I1(\u2.mem[27][7] ),
    .S(_04318_),
    .Z(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09302_ (.I(_04322_),
    .Z(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09303_ (.I(_04312_),
    .Z(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09304_ (.I0(_04269_),
    .I1(\u2.mem[27][8] ),
    .S(_04323_),
    .Z(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09305_ (.I(_04324_),
    .Z(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09306_ (.I0(_04272_),
    .I1(\u2.mem[27][9] ),
    .S(_04323_),
    .Z(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09307_ (.I(_04325_),
    .Z(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09308_ (.I0(_04274_),
    .I1(\u2.mem[27][10] ),
    .S(_04323_),
    .Z(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09309_ (.I(_04326_),
    .Z(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09310_ (.I0(_04276_),
    .I1(\u2.mem[27][11] ),
    .S(_04323_),
    .Z(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09311_ (.I(_04327_),
    .Z(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09312_ (.I(_04312_),
    .Z(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09313_ (.I0(_04278_),
    .I1(\u2.mem[27][12] ),
    .S(_04328_),
    .Z(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09314_ (.I(_04329_),
    .Z(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09315_ (.I0(_04281_),
    .I1(\u2.mem[27][13] ),
    .S(_04328_),
    .Z(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09316_ (.I(_04330_),
    .Z(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09317_ (.I0(_04283_),
    .I1(\u2.mem[27][14] ),
    .S(_04328_),
    .Z(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09318_ (.I(_04331_),
    .Z(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09319_ (.I0(_04285_),
    .I1(\u2.mem[27][15] ),
    .S(_04328_),
    .Z(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09320_ (.I(_04332_),
    .Z(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _09321_ (.A1(_03630_),
    .A2(_03540_),
    .A3(_03878_),
    .Z(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09322_ (.I(_04333_),
    .Z(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09323_ (.A1(_04011_),
    .A2(_04334_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09324_ (.I(_04335_),
    .Z(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09325_ (.I0(_04246_),
    .I1(\u2.mem[28][0] ),
    .S(_04336_),
    .Z(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09326_ (.I(_04337_),
    .Z(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09327_ (.I0(_04254_),
    .I1(\u2.mem[28][1] ),
    .S(_04336_),
    .Z(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09328_ (.I(_04338_),
    .Z(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09329_ (.I0(_04256_),
    .I1(\u2.mem[28][2] ),
    .S(_04336_),
    .Z(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09330_ (.I(_04339_),
    .Z(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09331_ (.I0(_04258_),
    .I1(\u2.mem[28][3] ),
    .S(_04336_),
    .Z(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09332_ (.I(_04340_),
    .Z(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09333_ (.I(_04335_),
    .Z(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09334_ (.I0(_04260_),
    .I1(\u2.mem[28][4] ),
    .S(_04341_),
    .Z(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09335_ (.I(_04342_),
    .Z(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09336_ (.I0(_04263_),
    .I1(\u2.mem[28][5] ),
    .S(_04341_),
    .Z(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09337_ (.I(_04343_),
    .Z(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09338_ (.I0(_04265_),
    .I1(\u2.mem[28][6] ),
    .S(_04341_),
    .Z(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09339_ (.I(_04344_),
    .Z(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09340_ (.I0(_04267_),
    .I1(\u2.mem[28][7] ),
    .S(_04341_),
    .Z(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09341_ (.I(_04345_),
    .Z(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09342_ (.I(_04335_),
    .Z(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09343_ (.I0(_04269_),
    .I1(\u2.mem[28][8] ),
    .S(_04346_),
    .Z(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09344_ (.I(_04347_),
    .Z(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09345_ (.I0(_04272_),
    .I1(\u2.mem[28][9] ),
    .S(_04346_),
    .Z(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09346_ (.I(_04348_),
    .Z(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09347_ (.I0(_04274_),
    .I1(\u2.mem[28][10] ),
    .S(_04346_),
    .Z(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09348_ (.I(_04349_),
    .Z(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09349_ (.I0(_04276_),
    .I1(\u2.mem[28][11] ),
    .S(_04346_),
    .Z(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09350_ (.I(_04350_),
    .Z(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09351_ (.I(_04335_),
    .Z(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09352_ (.I0(_04278_),
    .I1(\u2.mem[28][12] ),
    .S(_04351_),
    .Z(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09353_ (.I(_04352_),
    .Z(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09354_ (.I0(_04281_),
    .I1(\u2.mem[28][13] ),
    .S(_04351_),
    .Z(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09355_ (.I(_04353_),
    .Z(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09356_ (.I0(_04283_),
    .I1(\u2.mem[28][14] ),
    .S(_04351_),
    .Z(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09357_ (.I(_04354_),
    .Z(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09358_ (.I0(_04285_),
    .I1(\u2.mem[28][15] ),
    .S(_04351_),
    .Z(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09359_ (.I(_04355_),
    .Z(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09360_ (.I(_04118_),
    .Z(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09361_ (.A1(_03904_),
    .A2(_04250_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09362_ (.I(_04357_),
    .Z(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09363_ (.I0(_04356_),
    .I1(\u2.mem[29][0] ),
    .S(_04358_),
    .Z(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09364_ (.I(_04359_),
    .Z(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09365_ (.I(_04127_),
    .Z(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09366_ (.I0(_04360_),
    .I1(\u2.mem[29][1] ),
    .S(_04358_),
    .Z(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09367_ (.I(_04361_),
    .Z(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09368_ (.I(_04131_),
    .Z(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09369_ (.I0(_04362_),
    .I1(\u2.mem[29][2] ),
    .S(_04358_),
    .Z(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09370_ (.I(_04363_),
    .Z(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09371_ (.I(_04135_),
    .Z(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09372_ (.I0(_04364_),
    .I1(\u2.mem[29][3] ),
    .S(_04358_),
    .Z(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09373_ (.I(_04365_),
    .Z(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09374_ (.I(_04139_),
    .Z(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09375_ (.I(_04357_),
    .Z(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09376_ (.I0(_04366_),
    .I1(\u2.mem[29][4] ),
    .S(_04367_),
    .Z(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09377_ (.I(_04368_),
    .Z(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09378_ (.I(_04144_),
    .Z(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09379_ (.I0(_04369_),
    .I1(\u2.mem[29][5] ),
    .S(_04367_),
    .Z(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09380_ (.I(_04370_),
    .Z(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09381_ (.I(_04147_),
    .Z(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09382_ (.I0(_04371_),
    .I1(\u2.mem[29][6] ),
    .S(_04367_),
    .Z(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09383_ (.I(_04372_),
    .Z(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09384_ (.I(_04150_),
    .Z(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09385_ (.I0(_04373_),
    .I1(\u2.mem[29][7] ),
    .S(_04367_),
    .Z(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09386_ (.I(_04374_),
    .Z(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09387_ (.I(_04153_),
    .Z(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09388_ (.I(_04357_),
    .Z(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09389_ (.I0(_04375_),
    .I1(\u2.mem[29][8] ),
    .S(_04376_),
    .Z(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09390_ (.I(_04377_),
    .Z(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09391_ (.I(_04157_),
    .Z(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09392_ (.I0(_04378_),
    .I1(\u2.mem[29][9] ),
    .S(_04376_),
    .Z(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09393_ (.I(_04379_),
    .Z(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09394_ (.I(_04160_),
    .Z(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09395_ (.I0(_04380_),
    .I1(\u2.mem[29][10] ),
    .S(_04376_),
    .Z(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09396_ (.I(_04381_),
    .Z(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09397_ (.I(_04163_),
    .Z(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09398_ (.I0(_04382_),
    .I1(\u2.mem[29][11] ),
    .S(_04376_),
    .Z(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09399_ (.I(_04383_),
    .Z(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09400_ (.I(_04166_),
    .Z(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09401_ (.I(_04357_),
    .Z(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09402_ (.I0(_04384_),
    .I1(\u2.mem[29][12] ),
    .S(_04385_),
    .Z(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09403_ (.I(_04386_),
    .Z(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09404_ (.I(_04170_),
    .Z(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09405_ (.I0(_04387_),
    .I1(\u2.mem[29][13] ),
    .S(_04385_),
    .Z(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09406_ (.I(_04388_),
    .Z(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09407_ (.I(_04173_),
    .Z(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09408_ (.I0(_04389_),
    .I1(\u2.mem[29][14] ),
    .S(_04385_),
    .Z(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09409_ (.I(_04390_),
    .Z(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09410_ (.I(_04176_),
    .Z(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09411_ (.I0(_04391_),
    .I1(\u2.mem[29][15] ),
    .S(_04385_),
    .Z(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09412_ (.I(_04392_),
    .Z(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09413_ (.A1(_03581_),
    .A2(_03902_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09414_ (.I(_04393_),
    .Z(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09415_ (.A1(_04394_),
    .A2(_04011_),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09416_ (.I(_04395_),
    .Z(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09417_ (.I0(_04356_),
    .I1(\u2.mem[30][0] ),
    .S(_04396_),
    .Z(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09418_ (.I(_04397_),
    .Z(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09419_ (.I0(_04360_),
    .I1(\u2.mem[30][1] ),
    .S(_04396_),
    .Z(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09420_ (.I(_04398_),
    .Z(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09421_ (.I0(_04362_),
    .I1(\u2.mem[30][2] ),
    .S(_04396_),
    .Z(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09422_ (.I(_04399_),
    .Z(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09423_ (.I0(_04364_),
    .I1(\u2.mem[30][3] ),
    .S(_04396_),
    .Z(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09424_ (.I(_04400_),
    .Z(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09425_ (.I(_04395_),
    .Z(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09426_ (.I0(_04366_),
    .I1(\u2.mem[30][4] ),
    .S(_04401_),
    .Z(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09427_ (.I(_04402_),
    .Z(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09428_ (.I0(_04369_),
    .I1(\u2.mem[30][5] ),
    .S(_04401_),
    .Z(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09429_ (.I(_04403_),
    .Z(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09430_ (.I0(_04371_),
    .I1(\u2.mem[30][6] ),
    .S(_04401_),
    .Z(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09431_ (.I(_04404_),
    .Z(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09432_ (.I0(_04373_),
    .I1(\u2.mem[30][7] ),
    .S(_04401_),
    .Z(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09433_ (.I(_04405_),
    .Z(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09434_ (.I(_04395_),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09435_ (.I0(_04375_),
    .I1(\u2.mem[30][8] ),
    .S(_04406_),
    .Z(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09436_ (.I(_04407_),
    .Z(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09437_ (.I0(_04378_),
    .I1(\u2.mem[30][9] ),
    .S(_04406_),
    .Z(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09438_ (.I(_04408_),
    .Z(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09439_ (.I0(_04380_),
    .I1(\u2.mem[30][10] ),
    .S(_04406_),
    .Z(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09440_ (.I(_04409_),
    .Z(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09441_ (.I0(_04382_),
    .I1(\u2.mem[30][11] ),
    .S(_04406_),
    .Z(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09442_ (.I(_04410_),
    .Z(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09443_ (.I(_04395_),
    .Z(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09444_ (.I0(_04384_),
    .I1(\u2.mem[30][12] ),
    .S(_04411_),
    .Z(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09445_ (.I(_04412_),
    .Z(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09446_ (.I0(_04387_),
    .I1(\u2.mem[30][13] ),
    .S(_04411_),
    .Z(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09447_ (.I(_04413_),
    .Z(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09448_ (.I0(_04389_),
    .I1(\u2.mem[30][14] ),
    .S(_04411_),
    .Z(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09449_ (.I(_04414_),
    .Z(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09450_ (.I0(_04391_),
    .I1(\u2.mem[30][15] ),
    .S(_04411_),
    .Z(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09451_ (.I(_04415_),
    .Z(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09452_ (.A1(_03748_),
    .A2(_03902_),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09453_ (.I(_04416_),
    .Z(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09454_ (.A1(_04417_),
    .A2(_04011_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09455_ (.I(_04418_),
    .Z(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09456_ (.I0(_04356_),
    .I1(\u2.mem[31][0] ),
    .S(_04419_),
    .Z(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09457_ (.I(_04420_),
    .Z(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09458_ (.I0(_04360_),
    .I1(\u2.mem[31][1] ),
    .S(_04419_),
    .Z(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09459_ (.I(_04421_),
    .Z(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09460_ (.I0(_04362_),
    .I1(\u2.mem[31][2] ),
    .S(_04419_),
    .Z(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09461_ (.I(_04422_),
    .Z(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09462_ (.I0(_04364_),
    .I1(\u2.mem[31][3] ),
    .S(_04419_),
    .Z(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09463_ (.I(_04423_),
    .Z(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09464_ (.I(_04418_),
    .Z(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09465_ (.I0(_04366_),
    .I1(\u2.mem[31][4] ),
    .S(_04424_),
    .Z(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09466_ (.I(_04425_),
    .Z(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09467_ (.I0(_04369_),
    .I1(\u2.mem[31][5] ),
    .S(_04424_),
    .Z(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09468_ (.I(_04426_),
    .Z(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09469_ (.I0(_04371_),
    .I1(\u2.mem[31][6] ),
    .S(_04424_),
    .Z(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09470_ (.I(_04427_),
    .Z(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09471_ (.I0(_04373_),
    .I1(\u2.mem[31][7] ),
    .S(_04424_),
    .Z(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09472_ (.I(_04428_),
    .Z(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09473_ (.I(_04418_),
    .Z(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09474_ (.I0(_04375_),
    .I1(\u2.mem[31][8] ),
    .S(_04429_),
    .Z(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09475_ (.I(_04430_),
    .Z(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09476_ (.I0(_04378_),
    .I1(\u2.mem[31][9] ),
    .S(_04429_),
    .Z(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09477_ (.I(_04431_),
    .Z(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09478_ (.I0(_04380_),
    .I1(\u2.mem[31][10] ),
    .S(_04429_),
    .Z(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09479_ (.I(_04432_),
    .Z(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09480_ (.I0(_04382_),
    .I1(\u2.mem[31][11] ),
    .S(_04429_),
    .Z(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09481_ (.I(_04433_),
    .Z(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09482_ (.I(_04418_),
    .Z(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09483_ (.I0(_04384_),
    .I1(\u2.mem[31][12] ),
    .S(_04434_),
    .Z(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09484_ (.I(_04435_),
    .Z(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09485_ (.I0(_04387_),
    .I1(\u2.mem[31][13] ),
    .S(_04434_),
    .Z(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09486_ (.I(_04436_),
    .Z(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09487_ (.I0(_04389_),
    .I1(\u2.mem[31][14] ),
    .S(_04434_),
    .Z(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09488_ (.I(_04437_),
    .Z(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09489_ (.I0(_04391_),
    .I1(\u2.mem[31][15] ),
    .S(_04434_),
    .Z(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09490_ (.I(_04438_),
    .Z(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09491_ (.A1(_03984_),
    .A2(_03985_),
    .ZN(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09492_ (.A1(_03478_),
    .A2(_03986_),
    .A3(_04439_),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09493_ (.I(_04440_),
    .Z(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09494_ (.A1(_03983_),
    .A2(_04441_),
    .ZN(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09495_ (.I(_04442_),
    .Z(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09496_ (.I0(_04356_),
    .I1(\u2.mem[32][0] ),
    .S(_04443_),
    .Z(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09497_ (.I(_04444_),
    .Z(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09498_ (.I0(_04360_),
    .I1(\u2.mem[32][1] ),
    .S(_04443_),
    .Z(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09499_ (.I(_04445_),
    .Z(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09500_ (.I0(_04362_),
    .I1(\u2.mem[32][2] ),
    .S(_04443_),
    .Z(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09501_ (.I(_04446_),
    .Z(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09502_ (.I0(_04364_),
    .I1(\u2.mem[32][3] ),
    .S(_04443_),
    .Z(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09503_ (.I(_04447_),
    .Z(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09504_ (.I(_04442_),
    .Z(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09505_ (.I0(_04366_),
    .I1(\u2.mem[32][4] ),
    .S(_04448_),
    .Z(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09506_ (.I(_04449_),
    .Z(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09507_ (.I0(_04369_),
    .I1(\u2.mem[32][5] ),
    .S(_04448_),
    .Z(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09508_ (.I(_04450_),
    .Z(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09509_ (.I0(_04371_),
    .I1(\u2.mem[32][6] ),
    .S(_04448_),
    .Z(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09510_ (.I(_04451_),
    .Z(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09511_ (.I0(_04373_),
    .I1(\u2.mem[32][7] ),
    .S(_04448_),
    .Z(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09512_ (.I(_04452_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09513_ (.I(_04442_),
    .Z(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09514_ (.I0(_04375_),
    .I1(\u2.mem[32][8] ),
    .S(_04453_),
    .Z(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09515_ (.I(_04454_),
    .Z(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09516_ (.I0(_04378_),
    .I1(\u2.mem[32][9] ),
    .S(_04453_),
    .Z(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09517_ (.I(_04455_),
    .Z(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09518_ (.I0(_04380_),
    .I1(\u2.mem[32][10] ),
    .S(_04453_),
    .Z(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09519_ (.I(_04456_),
    .Z(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09520_ (.I0(_04382_),
    .I1(\u2.mem[32][11] ),
    .S(_04453_),
    .Z(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09521_ (.I(_04457_),
    .Z(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09522_ (.I(_04442_),
    .Z(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09523_ (.I0(_04384_),
    .I1(\u2.mem[32][12] ),
    .S(_04458_),
    .Z(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09524_ (.I(_04459_),
    .Z(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09525_ (.I0(_04387_),
    .I1(\u2.mem[32][13] ),
    .S(_04458_),
    .Z(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09526_ (.I(_04460_),
    .Z(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09527_ (.I0(_04389_),
    .I1(\u2.mem[32][14] ),
    .S(_04458_),
    .Z(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09528_ (.I(_04461_),
    .Z(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09529_ (.I0(_04391_),
    .I1(\u2.mem[32][15] ),
    .S(_04458_),
    .Z(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09530_ (.I(_04462_),
    .Z(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09531_ (.I(_04118_),
    .Z(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09532_ (.A1(_04013_),
    .A2(_04441_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09533_ (.I(_04464_),
    .Z(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09534_ (.I0(_04463_),
    .I1(\u2.mem[33][0] ),
    .S(_04465_),
    .Z(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09535_ (.I(_04466_),
    .Z(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09536_ (.I(_04127_),
    .Z(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09537_ (.I0(_04467_),
    .I1(\u2.mem[33][1] ),
    .S(_04465_),
    .Z(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09538_ (.I(_04468_),
    .Z(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09539_ (.I(_04131_),
    .Z(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09540_ (.I0(_04469_),
    .I1(\u2.mem[33][2] ),
    .S(_04465_),
    .Z(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09541_ (.I(_04470_),
    .Z(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09542_ (.I(_04135_),
    .Z(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09543_ (.I0(_04471_),
    .I1(\u2.mem[33][3] ),
    .S(_04465_),
    .Z(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09544_ (.I(_04472_),
    .Z(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09545_ (.I(_04139_),
    .Z(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09546_ (.I(_04464_),
    .Z(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09547_ (.I0(_04473_),
    .I1(\u2.mem[33][4] ),
    .S(_04474_),
    .Z(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09548_ (.I(_04475_),
    .Z(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09549_ (.I(_04144_),
    .Z(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09550_ (.I0(_04476_),
    .I1(\u2.mem[33][5] ),
    .S(_04474_),
    .Z(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09551_ (.I(_04477_),
    .Z(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09552_ (.I(_04147_),
    .Z(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09553_ (.I0(_04478_),
    .I1(\u2.mem[33][6] ),
    .S(_04474_),
    .Z(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09554_ (.I(_04479_),
    .Z(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09555_ (.I(_04150_),
    .Z(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09556_ (.I0(_04480_),
    .I1(\u2.mem[33][7] ),
    .S(_04474_),
    .Z(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09557_ (.I(_04481_),
    .Z(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09558_ (.I(_04153_),
    .Z(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09559_ (.I(_04464_),
    .Z(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09560_ (.I0(_04482_),
    .I1(\u2.mem[33][8] ),
    .S(_04483_),
    .Z(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09561_ (.I(_04484_),
    .Z(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09562_ (.I(_04157_),
    .Z(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09563_ (.I0(_04485_),
    .I1(\u2.mem[33][9] ),
    .S(_04483_),
    .Z(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09564_ (.I(_04486_),
    .Z(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09565_ (.I(_04160_),
    .Z(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09566_ (.I0(_04487_),
    .I1(\u2.mem[33][10] ),
    .S(_04483_),
    .Z(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09567_ (.I(_04488_),
    .Z(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09568_ (.I(_04163_),
    .Z(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09569_ (.I0(_04489_),
    .I1(\u2.mem[33][11] ),
    .S(_04483_),
    .Z(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09570_ (.I(_04490_),
    .Z(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09571_ (.I(_04166_),
    .Z(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09572_ (.I(_04464_),
    .Z(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09573_ (.I0(_04491_),
    .I1(\u2.mem[33][12] ),
    .S(_04492_),
    .Z(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09574_ (.I(_04493_),
    .Z(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09575_ (.I(_04170_),
    .Z(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09576_ (.I0(_04494_),
    .I1(\u2.mem[33][13] ),
    .S(_04492_),
    .Z(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09577_ (.I(_04495_),
    .Z(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09578_ (.I(_04173_),
    .Z(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09579_ (.I0(_04496_),
    .I1(\u2.mem[33][14] ),
    .S(_04492_),
    .Z(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09580_ (.I(_04497_),
    .Z(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09581_ (.I(_04176_),
    .Z(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09582_ (.I0(_04498_),
    .I1(\u2.mem[33][15] ),
    .S(_04492_),
    .Z(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09583_ (.I(_04499_),
    .Z(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09584_ (.A1(_03583_),
    .A2(_04441_),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09585_ (.I(_04500_),
    .Z(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09586_ (.I0(_04463_),
    .I1(\u2.mem[34][0] ),
    .S(_04501_),
    .Z(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09587_ (.I(_04502_),
    .Z(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09588_ (.I0(_04467_),
    .I1(\u2.mem[34][1] ),
    .S(_04501_),
    .Z(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09589_ (.I(_04503_),
    .Z(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09590_ (.I0(_04469_),
    .I1(\u2.mem[34][2] ),
    .S(_04501_),
    .Z(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09591_ (.I(_04504_),
    .Z(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09592_ (.I0(_04471_),
    .I1(\u2.mem[34][3] ),
    .S(_04501_),
    .Z(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09593_ (.I(_04505_),
    .Z(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09594_ (.I(_04500_),
    .Z(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09595_ (.I0(_04473_),
    .I1(\u2.mem[34][4] ),
    .S(_04506_),
    .Z(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09596_ (.I(_04507_),
    .Z(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09597_ (.I0(_04476_),
    .I1(\u2.mem[34][5] ),
    .S(_04506_),
    .Z(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09598_ (.I(_04508_),
    .Z(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09599_ (.I0(_04478_),
    .I1(\u2.mem[34][6] ),
    .S(_04506_),
    .Z(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09600_ (.I(_04509_),
    .Z(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09601_ (.I0(_04480_),
    .I1(\u2.mem[34][7] ),
    .S(_04506_),
    .Z(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09602_ (.I(_04510_),
    .Z(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09603_ (.I(_04500_),
    .Z(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09604_ (.I0(_04482_),
    .I1(\u2.mem[34][8] ),
    .S(_04511_),
    .Z(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09605_ (.I(_04512_),
    .Z(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09606_ (.I0(_04485_),
    .I1(\u2.mem[34][9] ),
    .S(_04511_),
    .Z(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09607_ (.I(_04513_),
    .Z(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09608_ (.I0(_04487_),
    .I1(\u2.mem[34][10] ),
    .S(_04511_),
    .Z(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09609_ (.I(_04514_),
    .Z(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09610_ (.I0(_04489_),
    .I1(\u2.mem[34][11] ),
    .S(_04511_),
    .Z(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09611_ (.I(_04515_),
    .Z(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09612_ (.I(_04500_),
    .Z(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09613_ (.I0(_04491_),
    .I1(\u2.mem[34][12] ),
    .S(_04516_),
    .Z(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09614_ (.I(_04517_),
    .Z(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09615_ (.I0(_04494_),
    .I1(\u2.mem[34][13] ),
    .S(_04516_),
    .Z(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09616_ (.I(_04518_),
    .Z(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09617_ (.I0(_04496_),
    .I1(\u2.mem[34][14] ),
    .S(_04516_),
    .Z(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09618_ (.I(_04519_),
    .Z(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09619_ (.I0(_04498_),
    .I1(\u2.mem[34][15] ),
    .S(_04516_),
    .Z(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09620_ (.I(_04520_),
    .Z(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09621_ (.A1(_04072_),
    .A2(_04441_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09622_ (.I(_04521_),
    .Z(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09623_ (.I0(_04463_),
    .I1(\u2.mem[35][0] ),
    .S(_04522_),
    .Z(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09624_ (.I(_04523_),
    .Z(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09625_ (.I0(_04467_),
    .I1(\u2.mem[35][1] ),
    .S(_04522_),
    .Z(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09626_ (.I(_04524_),
    .Z(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09627_ (.I0(_04469_),
    .I1(\u2.mem[35][2] ),
    .S(_04522_),
    .Z(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09628_ (.I(_04525_),
    .Z(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09629_ (.I0(_04471_),
    .I1(\u2.mem[35][3] ),
    .S(_04522_),
    .Z(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09630_ (.I(_04526_),
    .Z(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09631_ (.I(_04521_),
    .Z(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09632_ (.I0(_04473_),
    .I1(\u2.mem[35][4] ),
    .S(_04527_),
    .Z(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09633_ (.I(_04528_),
    .Z(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09634_ (.I0(_04476_),
    .I1(\u2.mem[35][5] ),
    .S(_04527_),
    .Z(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09635_ (.I(_04529_),
    .Z(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09636_ (.I0(_04478_),
    .I1(\u2.mem[35][6] ),
    .S(_04527_),
    .Z(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09637_ (.I(_04530_),
    .Z(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09638_ (.I0(_04480_),
    .I1(\u2.mem[35][7] ),
    .S(_04527_),
    .Z(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09639_ (.I(_04531_),
    .Z(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09640_ (.I(_04521_),
    .Z(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09641_ (.I0(_04482_),
    .I1(\u2.mem[35][8] ),
    .S(_04532_),
    .Z(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09642_ (.I(_04533_),
    .Z(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09643_ (.I0(_04485_),
    .I1(\u2.mem[35][9] ),
    .S(_04532_),
    .Z(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09644_ (.I(_04534_),
    .Z(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09645_ (.I0(_04487_),
    .I1(\u2.mem[35][10] ),
    .S(_04532_),
    .Z(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09646_ (.I(_04535_),
    .Z(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09647_ (.I0(_04489_),
    .I1(\u2.mem[35][11] ),
    .S(_04532_),
    .Z(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09648_ (.I(_04536_),
    .Z(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09649_ (.I(_04521_),
    .Z(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09650_ (.I0(_04491_),
    .I1(\u2.mem[35][12] ),
    .S(_04537_),
    .Z(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09651_ (.I(_04538_),
    .Z(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09652_ (.I0(_04494_),
    .I1(\u2.mem[35][13] ),
    .S(_04537_),
    .Z(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09653_ (.I(_04539_),
    .Z(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09654_ (.I0(_04496_),
    .I1(\u2.mem[35][14] ),
    .S(_04537_),
    .Z(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09655_ (.I(_04540_),
    .Z(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09656_ (.I0(_04498_),
    .I1(\u2.mem[35][15] ),
    .S(_04537_),
    .Z(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09657_ (.I(_04541_),
    .Z(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09658_ (.I(_04440_),
    .Z(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09659_ (.A1(_04095_),
    .A2(_04542_),
    .ZN(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09660_ (.I(_04543_),
    .Z(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09661_ (.I0(_04463_),
    .I1(\u2.mem[36][0] ),
    .S(_04544_),
    .Z(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09662_ (.I(_04545_),
    .Z(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09663_ (.I0(_04467_),
    .I1(\u2.mem[36][1] ),
    .S(_04544_),
    .Z(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09664_ (.I(_04546_),
    .Z(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09665_ (.I0(_04469_),
    .I1(\u2.mem[36][2] ),
    .S(_04544_),
    .Z(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09666_ (.I(_04547_),
    .Z(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09667_ (.I0(_04471_),
    .I1(\u2.mem[36][3] ),
    .S(_04544_),
    .Z(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09668_ (.I(_04548_),
    .Z(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09669_ (.I(_04543_),
    .Z(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09670_ (.I0(_04473_),
    .I1(\u2.mem[36][4] ),
    .S(_04549_),
    .Z(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09671_ (.I(_04550_),
    .Z(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09672_ (.I0(_04476_),
    .I1(\u2.mem[36][5] ),
    .S(_04549_),
    .Z(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09673_ (.I(_04551_),
    .Z(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09674_ (.I0(_04478_),
    .I1(\u2.mem[36][6] ),
    .S(_04549_),
    .Z(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09675_ (.I(_04552_),
    .Z(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09676_ (.I0(_04480_),
    .I1(\u2.mem[36][7] ),
    .S(_04549_),
    .Z(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09677_ (.I(_04553_),
    .Z(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09678_ (.I(_04543_),
    .Z(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09679_ (.I0(_04482_),
    .I1(\u2.mem[36][8] ),
    .S(_04554_),
    .Z(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09680_ (.I(_04555_),
    .Z(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09681_ (.I0(_04485_),
    .I1(\u2.mem[36][9] ),
    .S(_04554_),
    .Z(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09682_ (.I(_04556_),
    .Z(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09683_ (.I0(_04487_),
    .I1(\u2.mem[36][10] ),
    .S(_04554_),
    .Z(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09684_ (.I(_04557_),
    .Z(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09685_ (.I0(_04489_),
    .I1(\u2.mem[36][11] ),
    .S(_04554_),
    .Z(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09686_ (.I(_04558_),
    .Z(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09687_ (.I(_04543_),
    .Z(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09688_ (.I0(_04491_),
    .I1(\u2.mem[36][12] ),
    .S(_04559_),
    .Z(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09689_ (.I(_04560_),
    .Z(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09690_ (.I0(_04494_),
    .I1(\u2.mem[36][13] ),
    .S(_04559_),
    .Z(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09691_ (.I(_04561_),
    .Z(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09692_ (.I0(_04496_),
    .I1(\u2.mem[36][14] ),
    .S(_04559_),
    .Z(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09693_ (.I(_04562_),
    .Z(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09694_ (.I0(_04498_),
    .I1(\u2.mem[36][15] ),
    .S(_04559_),
    .Z(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09695_ (.I(_04563_),
    .Z(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09696_ (.I(_04117_),
    .Z(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09697_ (.I(_04564_),
    .Z(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09698_ (.A1(_04121_),
    .A2(_04542_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09699_ (.I(_04566_),
    .Z(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09700_ (.I0(_04565_),
    .I1(\u2.mem[37][0] ),
    .S(_04567_),
    .Z(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09701_ (.I(_04568_),
    .Z(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09702_ (.I(_04126_),
    .Z(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09703_ (.I(_04569_),
    .Z(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09704_ (.I0(_04570_),
    .I1(\u2.mem[37][1] ),
    .S(_04567_),
    .Z(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09705_ (.I(_04571_),
    .Z(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09706_ (.I(_04130_),
    .Z(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09707_ (.I(_04572_),
    .Z(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09708_ (.I0(_04573_),
    .I1(\u2.mem[37][2] ),
    .S(_04567_),
    .Z(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09709_ (.I(_04574_),
    .Z(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09710_ (.I(_04134_),
    .Z(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09711_ (.I(_04575_),
    .Z(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09712_ (.I0(_04576_),
    .I1(\u2.mem[37][3] ),
    .S(_04567_),
    .Z(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09713_ (.I(_04577_),
    .Z(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09714_ (.I(_04138_),
    .Z(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09715_ (.I(_04578_),
    .Z(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09716_ (.I(_04566_),
    .Z(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09717_ (.I0(_04579_),
    .I1(\u2.mem[37][4] ),
    .S(_04580_),
    .Z(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09718_ (.I(_04581_),
    .Z(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09719_ (.I(_04143_),
    .Z(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09720_ (.I(_04582_),
    .Z(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09721_ (.I0(_04583_),
    .I1(\u2.mem[37][5] ),
    .S(_04580_),
    .Z(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09722_ (.I(_04584_),
    .Z(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09723_ (.I(\data_in_trans[6].data_sync ),
    .Z(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09724_ (.I(_04585_),
    .Z(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09725_ (.I0(_04586_),
    .I1(\u2.mem[37][6] ),
    .S(_04580_),
    .Z(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09726_ (.I(_04587_),
    .Z(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09727_ (.I(\data_in_trans[7].data_sync ),
    .Z(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09728_ (.I(_04588_),
    .Z(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09729_ (.I0(_04589_),
    .I1(\u2.mem[37][7] ),
    .S(_04580_),
    .Z(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09730_ (.I(_04590_),
    .Z(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09731_ (.I(\data_in_trans[8].data_sync ),
    .Z(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09732_ (.I(_04591_),
    .Z(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09733_ (.I(_04566_),
    .Z(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09734_ (.I0(_04592_),
    .I1(\u2.mem[37][8] ),
    .S(_04593_),
    .Z(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09735_ (.I(_04594_),
    .Z(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09736_ (.I(\data_in_trans[9].data_sync ),
    .Z(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09737_ (.I(_04595_),
    .Z(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09738_ (.I0(_04596_),
    .I1(\u2.mem[37][9] ),
    .S(_04593_),
    .Z(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09739_ (.I(_04597_),
    .Z(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09740_ (.I(\data_in_trans[10].data_sync ),
    .Z(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09741_ (.I(_04598_),
    .Z(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09742_ (.I0(_04599_),
    .I1(\u2.mem[37][10] ),
    .S(_04593_),
    .Z(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09743_ (.I(_04600_),
    .Z(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09744_ (.I(\data_in_trans[11].data_sync ),
    .Z(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09745_ (.I(_04601_),
    .Z(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09746_ (.I0(_04602_),
    .I1(\u2.mem[37][11] ),
    .S(_04593_),
    .Z(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09747_ (.I(_04603_),
    .Z(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09748_ (.I(\data_in_trans[12].data_sync ),
    .Z(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09749_ (.I(_04604_),
    .Z(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09750_ (.I(_04566_),
    .Z(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09751_ (.I0(_04605_),
    .I1(\u2.mem[37][12] ),
    .S(_04606_),
    .Z(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09752_ (.I(_04607_),
    .Z(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09753_ (.I(\data_in_trans[13].data_sync ),
    .Z(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09754_ (.I(_04608_),
    .Z(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09755_ (.I0(_04609_),
    .I1(\u2.mem[37][13] ),
    .S(_04606_),
    .Z(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09756_ (.I(_04610_),
    .Z(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09757_ (.I(\data_in_trans[14].data_sync ),
    .Z(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09758_ (.I(_04611_),
    .Z(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09759_ (.I0(_04612_),
    .I1(\u2.mem[37][14] ),
    .S(_04606_),
    .Z(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09760_ (.I(_04613_),
    .Z(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09761_ (.I(\data_in_trans[15].data_sync ),
    .Z(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09762_ (.I(_04614_),
    .Z(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09763_ (.I0(_04615_),
    .I1(\u2.mem[37][15] ),
    .S(_04606_),
    .Z(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09764_ (.I(_04616_),
    .Z(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09765_ (.A1(_04180_),
    .A2(_04542_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09766_ (.I(_04617_),
    .Z(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09767_ (.I0(_04565_),
    .I1(\u2.mem[38][0] ),
    .S(_04618_),
    .Z(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09768_ (.I(_04619_),
    .Z(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09769_ (.I0(_04570_),
    .I1(\u2.mem[38][1] ),
    .S(_04618_),
    .Z(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09770_ (.I(_04620_),
    .Z(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09771_ (.I0(_04573_),
    .I1(\u2.mem[38][2] ),
    .S(_04618_),
    .Z(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09772_ (.I(_04621_),
    .Z(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09773_ (.I0(_04576_),
    .I1(\u2.mem[38][3] ),
    .S(_04618_),
    .Z(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09774_ (.I(_04622_),
    .Z(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09775_ (.I(_04617_),
    .Z(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09776_ (.I0(_04579_),
    .I1(\u2.mem[38][4] ),
    .S(_04623_),
    .Z(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09777_ (.I(_04624_),
    .Z(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09778_ (.I0(_04583_),
    .I1(\u2.mem[38][5] ),
    .S(_04623_),
    .Z(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09779_ (.I(_04625_),
    .Z(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09780_ (.I0(_04586_),
    .I1(\u2.mem[38][6] ),
    .S(_04623_),
    .Z(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09781_ (.I(_04626_),
    .Z(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09782_ (.I0(_04589_),
    .I1(\u2.mem[38][7] ),
    .S(_04623_),
    .Z(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09783_ (.I(_04627_),
    .Z(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09784_ (.I(_04617_),
    .Z(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09785_ (.I0(_04592_),
    .I1(\u2.mem[38][8] ),
    .S(_04628_),
    .Z(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09786_ (.I(_04629_),
    .Z(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09787_ (.I0(_04596_),
    .I1(\u2.mem[38][9] ),
    .S(_04628_),
    .Z(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09788_ (.I(_04630_),
    .Z(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09789_ (.I0(_04599_),
    .I1(\u2.mem[38][10] ),
    .S(_04628_),
    .Z(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09790_ (.I(_04631_),
    .Z(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09791_ (.I0(_04602_),
    .I1(\u2.mem[38][11] ),
    .S(_04628_),
    .Z(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09792_ (.I(_04632_),
    .Z(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09793_ (.I(_04617_),
    .Z(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09794_ (.I0(_04605_),
    .I1(\u2.mem[38][12] ),
    .S(_04633_),
    .Z(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09795_ (.I(_04634_),
    .Z(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09796_ (.I0(_04609_),
    .I1(\u2.mem[38][13] ),
    .S(_04633_),
    .Z(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09797_ (.I(_04635_),
    .Z(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09798_ (.I0(_04612_),
    .I1(\u2.mem[38][14] ),
    .S(_04633_),
    .Z(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09799_ (.I(_04636_),
    .Z(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09800_ (.I0(_04615_),
    .I1(\u2.mem[38][15] ),
    .S(_04633_),
    .Z(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09801_ (.I(_04637_),
    .Z(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09802_ (.A1(_03752_),
    .A2(_04542_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09803_ (.I(_04638_),
    .Z(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09804_ (.I0(_04565_),
    .I1(\u2.mem[39][0] ),
    .S(_04639_),
    .Z(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09805_ (.I(_04640_),
    .Z(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09806_ (.I0(_04570_),
    .I1(\u2.mem[39][1] ),
    .S(_04639_),
    .Z(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09807_ (.I(_04641_),
    .Z(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09808_ (.I0(_04573_),
    .I1(\u2.mem[39][2] ),
    .S(_04639_),
    .Z(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09809_ (.I(_04642_),
    .Z(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09810_ (.I0(_04576_),
    .I1(\u2.mem[39][3] ),
    .S(_04639_),
    .Z(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09811_ (.I(_04643_),
    .Z(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09812_ (.I(_04638_),
    .Z(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09813_ (.I0(_04579_),
    .I1(\u2.mem[39][4] ),
    .S(_04644_),
    .Z(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09814_ (.I(_04645_),
    .Z(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09815_ (.I0(_04583_),
    .I1(\u2.mem[39][5] ),
    .S(_04644_),
    .Z(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09816_ (.I(_04646_),
    .Z(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09817_ (.I0(_04586_),
    .I1(\u2.mem[39][6] ),
    .S(_04644_),
    .Z(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09818_ (.I(_04647_),
    .Z(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09819_ (.I0(_04589_),
    .I1(\u2.mem[39][7] ),
    .S(_04644_),
    .Z(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09820_ (.I(_04648_),
    .Z(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09821_ (.I(_04638_),
    .Z(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09822_ (.I0(_04592_),
    .I1(\u2.mem[39][8] ),
    .S(_04649_),
    .Z(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09823_ (.I(_04650_),
    .Z(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09824_ (.I0(_04596_),
    .I1(\u2.mem[39][9] ),
    .S(_04649_),
    .Z(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09825_ (.I(_04651_),
    .Z(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09826_ (.I0(_04599_),
    .I1(\u2.mem[39][10] ),
    .S(_04649_),
    .Z(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09827_ (.I(_04652_),
    .Z(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09828_ (.I0(_04602_),
    .I1(\u2.mem[39][11] ),
    .S(_04649_),
    .Z(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09829_ (.I(_04653_),
    .Z(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09830_ (.I(_04638_),
    .Z(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09831_ (.I0(_04605_),
    .I1(\u2.mem[39][12] ),
    .S(_04654_),
    .Z(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09832_ (.I(_04655_),
    .Z(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09833_ (.I0(_04609_),
    .I1(\u2.mem[39][13] ),
    .S(_04654_),
    .Z(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09834_ (.I(_04656_),
    .Z(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09835_ (.I0(_04612_),
    .I1(\u2.mem[39][14] ),
    .S(_04654_),
    .Z(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09836_ (.I(_04657_),
    .Z(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09837_ (.I0(_04615_),
    .I1(\u2.mem[39][15] ),
    .S(_04654_),
    .Z(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09838_ (.I(_04658_),
    .Z(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09839_ (.I(_04440_),
    .Z(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09840_ (.A1(_04224_),
    .A2(_04659_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09841_ (.I(_04660_),
    .Z(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09842_ (.I0(_04565_),
    .I1(\u2.mem[40][0] ),
    .S(_04661_),
    .Z(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09843_ (.I(_04662_),
    .Z(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09844_ (.I0(_04570_),
    .I1(\u2.mem[40][1] ),
    .S(_04661_),
    .Z(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09845_ (.I(_04663_),
    .Z(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09846_ (.I0(_04573_),
    .I1(\u2.mem[40][2] ),
    .S(_04661_),
    .Z(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09847_ (.I(_04664_),
    .Z(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09848_ (.I0(_04576_),
    .I1(\u2.mem[40][3] ),
    .S(_04661_),
    .Z(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09849_ (.I(_04665_),
    .Z(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09850_ (.I(_04660_),
    .Z(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09851_ (.I0(_04579_),
    .I1(\u2.mem[40][4] ),
    .S(_04666_),
    .Z(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09852_ (.I(_04667_),
    .Z(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09853_ (.I0(_04583_),
    .I1(\u2.mem[40][5] ),
    .S(_04666_),
    .Z(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09854_ (.I(_04668_),
    .Z(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09855_ (.I0(_04586_),
    .I1(\u2.mem[40][6] ),
    .S(_04666_),
    .Z(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09856_ (.I(_04669_),
    .Z(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09857_ (.I0(_04589_),
    .I1(\u2.mem[40][7] ),
    .S(_04666_),
    .Z(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09858_ (.I(_04670_),
    .Z(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09859_ (.I(_04660_),
    .Z(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09860_ (.I0(_04592_),
    .I1(\u2.mem[40][8] ),
    .S(_04671_),
    .Z(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09861_ (.I(_04672_),
    .Z(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09862_ (.I0(_04596_),
    .I1(\u2.mem[40][9] ),
    .S(_04671_),
    .Z(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09863_ (.I(_04673_),
    .Z(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09864_ (.I0(_04599_),
    .I1(\u2.mem[40][10] ),
    .S(_04671_),
    .Z(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09865_ (.I(_04674_),
    .Z(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09866_ (.I0(_04602_),
    .I1(\u2.mem[40][11] ),
    .S(_04671_),
    .Z(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09867_ (.I(_04675_),
    .Z(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09868_ (.I(_04660_),
    .Z(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09869_ (.I0(_04605_),
    .I1(\u2.mem[40][12] ),
    .S(_04676_),
    .Z(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09870_ (.I(_04677_),
    .Z(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09871_ (.I0(_04609_),
    .I1(\u2.mem[40][13] ),
    .S(_04676_),
    .Z(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09872_ (.I(_04678_),
    .Z(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09873_ (.I0(_04612_),
    .I1(\u2.mem[40][14] ),
    .S(_04676_),
    .Z(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09874_ (.I(_04679_),
    .Z(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09875_ (.I0(_04615_),
    .I1(\u2.mem[40][15] ),
    .S(_04676_),
    .Z(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09876_ (.I(_04680_),
    .Z(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09877_ (.I(_04564_),
    .Z(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09878_ (.A1(_04249_),
    .A2(_04659_),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09879_ (.I(_04682_),
    .Z(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09880_ (.I0(_04681_),
    .I1(\u2.mem[41][0] ),
    .S(_04683_),
    .Z(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09881_ (.I(_04684_),
    .Z(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09882_ (.I(_04569_),
    .Z(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09883_ (.I0(_04685_),
    .I1(\u2.mem[41][1] ),
    .S(_04683_),
    .Z(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09884_ (.I(_04686_),
    .Z(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09885_ (.I(_04572_),
    .Z(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09886_ (.I0(_04687_),
    .I1(\u2.mem[41][2] ),
    .S(_04683_),
    .Z(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09887_ (.I(_04688_),
    .Z(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09888_ (.I(_04575_),
    .Z(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09889_ (.I0(_04689_),
    .I1(\u2.mem[41][3] ),
    .S(_04683_),
    .Z(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09890_ (.I(_04690_),
    .Z(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09891_ (.I(_04578_),
    .Z(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09892_ (.I(_04682_),
    .Z(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09893_ (.I0(_04691_),
    .I1(\u2.mem[41][4] ),
    .S(_04692_),
    .Z(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09894_ (.I(_04693_),
    .Z(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09895_ (.I(_04582_),
    .Z(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09896_ (.I0(_04694_),
    .I1(\u2.mem[41][5] ),
    .S(_04692_),
    .Z(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09897_ (.I(_04695_),
    .Z(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09898_ (.I(_04585_),
    .Z(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09899_ (.I0(_04696_),
    .I1(\u2.mem[41][6] ),
    .S(_04692_),
    .Z(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09900_ (.I(_04697_),
    .Z(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09901_ (.I(_04588_),
    .Z(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09902_ (.I0(_04698_),
    .I1(\u2.mem[41][7] ),
    .S(_04692_),
    .Z(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09903_ (.I(_04699_),
    .Z(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09904_ (.I(_04591_),
    .Z(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09905_ (.I(_04682_),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09906_ (.I0(_04700_),
    .I1(\u2.mem[41][8] ),
    .S(_04701_),
    .Z(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09907_ (.I(_04702_),
    .Z(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09908_ (.I(_04595_),
    .Z(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09909_ (.I0(_04703_),
    .I1(\u2.mem[41][9] ),
    .S(_04701_),
    .Z(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09910_ (.I(_04704_),
    .Z(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09911_ (.I(_04598_),
    .Z(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09912_ (.I0(_04705_),
    .I1(\u2.mem[41][10] ),
    .S(_04701_),
    .Z(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09913_ (.I(_04706_),
    .Z(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09914_ (.I(_04601_),
    .Z(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09915_ (.I0(_04707_),
    .I1(\u2.mem[41][11] ),
    .S(_04701_),
    .Z(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09916_ (.I(_04708_),
    .Z(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09917_ (.I(_04604_),
    .Z(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09918_ (.I(_04682_),
    .Z(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09919_ (.I0(_04709_),
    .I1(\u2.mem[41][12] ),
    .S(_04710_),
    .Z(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09920_ (.I(_04711_),
    .Z(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09921_ (.I(_04608_),
    .Z(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09922_ (.I0(_04712_),
    .I1(\u2.mem[41][13] ),
    .S(_04710_),
    .Z(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09923_ (.I(_04713_),
    .Z(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09924_ (.I(_04611_),
    .Z(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09925_ (.I0(_04714_),
    .I1(\u2.mem[41][14] ),
    .S(_04710_),
    .Z(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09926_ (.I(_04715_),
    .Z(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09927_ (.I(_04614_),
    .Z(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09928_ (.I0(_04716_),
    .I1(\u2.mem[41][15] ),
    .S(_04710_),
    .Z(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09929_ (.I(_04717_),
    .Z(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09930_ (.A1(_04288_),
    .A2(_04659_),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09931_ (.I(_04718_),
    .Z(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09932_ (.I0(_04681_),
    .I1(\u2.mem[42][0] ),
    .S(_04719_),
    .Z(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09933_ (.I(_04720_),
    .Z(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09934_ (.I0(_04685_),
    .I1(\u2.mem[42][1] ),
    .S(_04719_),
    .Z(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09935_ (.I(_04721_),
    .Z(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09936_ (.I0(_04687_),
    .I1(\u2.mem[42][2] ),
    .S(_04719_),
    .Z(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09937_ (.I(_04722_),
    .Z(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09938_ (.I0(_04689_),
    .I1(\u2.mem[42][3] ),
    .S(_04719_),
    .Z(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09939_ (.I(_04723_),
    .Z(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09940_ (.I(_04718_),
    .Z(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09941_ (.I0(_04691_),
    .I1(\u2.mem[42][4] ),
    .S(_04724_),
    .Z(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09942_ (.I(_04725_),
    .Z(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09943_ (.I0(_04694_),
    .I1(\u2.mem[42][5] ),
    .S(_04724_),
    .Z(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09944_ (.I(_04726_),
    .Z(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09945_ (.I0(_04696_),
    .I1(\u2.mem[42][6] ),
    .S(_04724_),
    .Z(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09946_ (.I(_04727_),
    .Z(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09947_ (.I0(_04698_),
    .I1(\u2.mem[42][7] ),
    .S(_04724_),
    .Z(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09948_ (.I(_04728_),
    .Z(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09949_ (.I(_04718_),
    .Z(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09950_ (.I0(_04700_),
    .I1(\u2.mem[42][8] ),
    .S(_04729_),
    .Z(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09951_ (.I(_04730_),
    .Z(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09952_ (.I0(_04703_),
    .I1(\u2.mem[42][9] ),
    .S(_04729_),
    .Z(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09953_ (.I(_04731_),
    .Z(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09954_ (.I0(_04705_),
    .I1(\u2.mem[42][10] ),
    .S(_04729_),
    .Z(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09955_ (.I(_04732_),
    .Z(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09956_ (.I0(_04707_),
    .I1(\u2.mem[42][11] ),
    .S(_04729_),
    .Z(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09957_ (.I(_04733_),
    .Z(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09958_ (.I(_04718_),
    .Z(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09959_ (.I0(_04709_),
    .I1(\u2.mem[42][12] ),
    .S(_04734_),
    .Z(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09960_ (.I(_04735_),
    .Z(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09961_ (.I0(_04712_),
    .I1(\u2.mem[42][13] ),
    .S(_04734_),
    .Z(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09962_ (.I(_04736_),
    .Z(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09963_ (.I0(_04714_),
    .I1(\u2.mem[42][14] ),
    .S(_04734_),
    .Z(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09964_ (.I(_04737_),
    .Z(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09965_ (.I0(_04716_),
    .I1(\u2.mem[42][15] ),
    .S(_04734_),
    .Z(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09966_ (.I(_04738_),
    .Z(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09967_ (.A1(_04311_),
    .A2(_04659_),
    .ZN(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09968_ (.I(_04739_),
    .Z(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09969_ (.I0(_04681_),
    .I1(\u2.mem[43][0] ),
    .S(_04740_),
    .Z(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09970_ (.I(_04741_),
    .Z(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09971_ (.I0(_04685_),
    .I1(\u2.mem[43][1] ),
    .S(_04740_),
    .Z(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09972_ (.I(_04742_),
    .Z(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09973_ (.I0(_04687_),
    .I1(\u2.mem[43][2] ),
    .S(_04740_),
    .Z(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09974_ (.I(_04743_),
    .Z(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09975_ (.I0(_04689_),
    .I1(\u2.mem[43][3] ),
    .S(_04740_),
    .Z(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09976_ (.I(_04744_),
    .Z(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09977_ (.I(_04739_),
    .Z(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09978_ (.I0(_04691_),
    .I1(\u2.mem[43][4] ),
    .S(_04745_),
    .Z(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09979_ (.I(_04746_),
    .Z(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09980_ (.I0(_04694_),
    .I1(\u2.mem[43][5] ),
    .S(_04745_),
    .Z(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09981_ (.I(_04747_),
    .Z(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09982_ (.I0(_04696_),
    .I1(\u2.mem[43][6] ),
    .S(_04745_),
    .Z(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09983_ (.I(_04748_),
    .Z(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09984_ (.I0(_04698_),
    .I1(\u2.mem[43][7] ),
    .S(_04745_),
    .Z(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09985_ (.I(_04749_),
    .Z(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09986_ (.I(_04739_),
    .Z(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09987_ (.I0(_04700_),
    .I1(\u2.mem[43][8] ),
    .S(_04750_),
    .Z(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09988_ (.I(_04751_),
    .Z(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09989_ (.I0(_04703_),
    .I1(\u2.mem[43][9] ),
    .S(_04750_),
    .Z(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09990_ (.I(_04752_),
    .Z(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09991_ (.I0(_04705_),
    .I1(\u2.mem[43][10] ),
    .S(_04750_),
    .Z(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09992_ (.I(_04753_),
    .Z(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09993_ (.I0(_04707_),
    .I1(\u2.mem[43][11] ),
    .S(_04750_),
    .Z(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09994_ (.I(_04754_),
    .Z(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09995_ (.I(_04739_),
    .Z(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09996_ (.I0(_04709_),
    .I1(\u2.mem[43][12] ),
    .S(_04755_),
    .Z(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09997_ (.I(_04756_),
    .Z(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09998_ (.I0(_04712_),
    .I1(\u2.mem[43][13] ),
    .S(_04755_),
    .Z(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09999_ (.I(_04757_),
    .Z(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10000_ (.I0(_04714_),
    .I1(\u2.mem[43][14] ),
    .S(_04755_),
    .Z(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10001_ (.I(_04758_),
    .Z(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10002_ (.I0(_04716_),
    .I1(\u2.mem[43][15] ),
    .S(_04755_),
    .Z(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10003_ (.I(_04759_),
    .Z(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10004_ (.I(_04440_),
    .Z(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10005_ (.A1(_04334_),
    .A2(_04760_),
    .ZN(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10006_ (.I(_04761_),
    .Z(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10007_ (.I0(_04681_),
    .I1(\u2.mem[44][0] ),
    .S(_04762_),
    .Z(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10008_ (.I(_04763_),
    .Z(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10009_ (.I0(_04685_),
    .I1(\u2.mem[44][1] ),
    .S(_04762_),
    .Z(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10010_ (.I(_04764_),
    .Z(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10011_ (.I0(_04687_),
    .I1(\u2.mem[44][2] ),
    .S(_04762_),
    .Z(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10012_ (.I(_04765_),
    .Z(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10013_ (.I0(_04689_),
    .I1(\u2.mem[44][3] ),
    .S(_04762_),
    .Z(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10014_ (.I(_04766_),
    .Z(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10015_ (.I(_04761_),
    .Z(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10016_ (.I0(_04691_),
    .I1(\u2.mem[44][4] ),
    .S(_04767_),
    .Z(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10017_ (.I(_04768_),
    .Z(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10018_ (.I0(_04694_),
    .I1(\u2.mem[44][5] ),
    .S(_04767_),
    .Z(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10019_ (.I(_04769_),
    .Z(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10020_ (.I0(_04696_),
    .I1(\u2.mem[44][6] ),
    .S(_04767_),
    .Z(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10021_ (.I(_04770_),
    .Z(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10022_ (.I0(_04698_),
    .I1(\u2.mem[44][7] ),
    .S(_04767_),
    .Z(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10023_ (.I(_04771_),
    .Z(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10024_ (.I(_04761_),
    .Z(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10025_ (.I0(_04700_),
    .I1(\u2.mem[44][8] ),
    .S(_04772_),
    .Z(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10026_ (.I(_04773_),
    .Z(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10027_ (.I0(_04703_),
    .I1(\u2.mem[44][9] ),
    .S(_04772_),
    .Z(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10028_ (.I(_04774_),
    .Z(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10029_ (.I0(_04705_),
    .I1(\u2.mem[44][10] ),
    .S(_04772_),
    .Z(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10030_ (.I(_04775_),
    .Z(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10031_ (.I0(_04707_),
    .I1(\u2.mem[44][11] ),
    .S(_04772_),
    .Z(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10032_ (.I(_04776_),
    .Z(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10033_ (.I(_04761_),
    .Z(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10034_ (.I0(_04709_),
    .I1(\u2.mem[44][12] ),
    .S(_04777_),
    .Z(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10035_ (.I(_04778_),
    .Z(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10036_ (.I0(_04712_),
    .I1(\u2.mem[44][13] ),
    .S(_04777_),
    .Z(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10037_ (.I(_04779_),
    .Z(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10038_ (.I0(_04714_),
    .I1(\u2.mem[44][14] ),
    .S(_04777_),
    .Z(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10039_ (.I(_04780_),
    .Z(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10040_ (.I0(_04716_),
    .I1(\u2.mem[44][15] ),
    .S(_04777_),
    .Z(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10041_ (.I(_04781_),
    .Z(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10042_ (.I(_04564_),
    .Z(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10043_ (.A1(_03904_),
    .A2(_04760_),
    .ZN(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10044_ (.I(_04783_),
    .Z(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10045_ (.I0(_04782_),
    .I1(\u2.mem[45][0] ),
    .S(_04784_),
    .Z(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10046_ (.I(_04785_),
    .Z(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10047_ (.I(_04569_),
    .Z(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10048_ (.I0(_04786_),
    .I1(\u2.mem[45][1] ),
    .S(_04784_),
    .Z(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10049_ (.I(_04787_),
    .Z(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10050_ (.I(_04572_),
    .Z(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10051_ (.I0(_04788_),
    .I1(\u2.mem[45][2] ),
    .S(_04784_),
    .Z(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10052_ (.I(_04789_),
    .Z(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10053_ (.I(_04575_),
    .Z(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10054_ (.I0(_04790_),
    .I1(\u2.mem[45][3] ),
    .S(_04784_),
    .Z(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10055_ (.I(_04791_),
    .Z(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10056_ (.I(_04578_),
    .Z(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10057_ (.I(_04783_),
    .Z(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10058_ (.I0(_04792_),
    .I1(\u2.mem[45][4] ),
    .S(_04793_),
    .Z(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10059_ (.I(_04794_),
    .Z(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10060_ (.I(_04582_),
    .Z(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10061_ (.I0(_04795_),
    .I1(\u2.mem[45][5] ),
    .S(_04793_),
    .Z(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10062_ (.I(_04796_),
    .Z(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10063_ (.I(_04585_),
    .Z(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10064_ (.I0(_04797_),
    .I1(\u2.mem[45][6] ),
    .S(_04793_),
    .Z(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10065_ (.I(_04798_),
    .Z(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10066_ (.I(_04588_),
    .Z(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10067_ (.I0(_04799_),
    .I1(\u2.mem[45][7] ),
    .S(_04793_),
    .Z(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10068_ (.I(_04800_),
    .Z(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10069_ (.I(_04591_),
    .Z(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10070_ (.I(_04783_),
    .Z(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10071_ (.I0(_04801_),
    .I1(\u2.mem[45][8] ),
    .S(_04802_),
    .Z(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10072_ (.I(_04803_),
    .Z(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10073_ (.I(_04595_),
    .Z(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10074_ (.I0(_04804_),
    .I1(\u2.mem[45][9] ),
    .S(_04802_),
    .Z(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10075_ (.I(_04805_),
    .Z(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10076_ (.I(_04598_),
    .Z(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10077_ (.I0(_04806_),
    .I1(\u2.mem[45][10] ),
    .S(_04802_),
    .Z(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10078_ (.I(_04807_),
    .Z(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10079_ (.I(_04601_),
    .Z(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10080_ (.I0(_04808_),
    .I1(\u2.mem[45][11] ),
    .S(_04802_),
    .Z(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10081_ (.I(_04809_),
    .Z(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10082_ (.I(_04604_),
    .Z(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10083_ (.I(_04783_),
    .Z(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10084_ (.I0(_04810_),
    .I1(\u2.mem[45][12] ),
    .S(_04811_),
    .Z(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10085_ (.I(_04812_),
    .Z(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10086_ (.I(_04608_),
    .Z(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10087_ (.I0(_04813_),
    .I1(\u2.mem[45][13] ),
    .S(_04811_),
    .Z(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10088_ (.I(_04814_),
    .Z(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10089_ (.I(_04611_),
    .Z(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10090_ (.I0(_04815_),
    .I1(\u2.mem[45][14] ),
    .S(_04811_),
    .Z(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10091_ (.I(_04816_),
    .Z(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10092_ (.I(_04614_),
    .Z(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10093_ (.I0(_04817_),
    .I1(\u2.mem[45][15] ),
    .S(_04811_),
    .Z(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10094_ (.I(_04818_),
    .Z(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10095_ (.A1(_04394_),
    .A2(_04760_),
    .ZN(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10096_ (.I(_04819_),
    .Z(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10097_ (.I0(_04782_),
    .I1(\u2.mem[46][0] ),
    .S(_04820_),
    .Z(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10098_ (.I(_04821_),
    .Z(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10099_ (.I0(_04786_),
    .I1(\u2.mem[46][1] ),
    .S(_04820_),
    .Z(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10100_ (.I(_04822_),
    .Z(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10101_ (.I0(_04788_),
    .I1(\u2.mem[46][2] ),
    .S(_04820_),
    .Z(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10102_ (.I(_04823_),
    .Z(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10103_ (.I0(_04790_),
    .I1(\u2.mem[46][3] ),
    .S(_04820_),
    .Z(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10104_ (.I(_04824_),
    .Z(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10105_ (.I(_04819_),
    .Z(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10106_ (.I0(_04792_),
    .I1(\u2.mem[46][4] ),
    .S(_04825_),
    .Z(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10107_ (.I(_04826_),
    .Z(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10108_ (.I0(_04795_),
    .I1(\u2.mem[46][5] ),
    .S(_04825_),
    .Z(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10109_ (.I(_04827_),
    .Z(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10110_ (.I0(_04797_),
    .I1(\u2.mem[46][6] ),
    .S(_04825_),
    .Z(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10111_ (.I(_04828_),
    .Z(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10112_ (.I0(_04799_),
    .I1(\u2.mem[46][7] ),
    .S(_04825_),
    .Z(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10113_ (.I(_04829_),
    .Z(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10114_ (.I(_04819_),
    .Z(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10115_ (.I0(_04801_),
    .I1(\u2.mem[46][8] ),
    .S(_04830_),
    .Z(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10116_ (.I(_04831_),
    .Z(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10117_ (.I0(_04804_),
    .I1(\u2.mem[46][9] ),
    .S(_04830_),
    .Z(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10118_ (.I(_04832_),
    .Z(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10119_ (.I0(_04806_),
    .I1(\u2.mem[46][10] ),
    .S(_04830_),
    .Z(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10120_ (.I(_04833_),
    .Z(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10121_ (.I0(_04808_),
    .I1(\u2.mem[46][11] ),
    .S(_04830_),
    .Z(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10122_ (.I(_04834_),
    .Z(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10123_ (.I(_04819_),
    .Z(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10124_ (.I0(_04810_),
    .I1(\u2.mem[46][12] ),
    .S(_04835_),
    .Z(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10125_ (.I(_04836_),
    .Z(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10126_ (.I0(_04813_),
    .I1(\u2.mem[46][13] ),
    .S(_04835_),
    .Z(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10127_ (.I(_04837_),
    .Z(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10128_ (.I0(_04815_),
    .I1(\u2.mem[46][14] ),
    .S(_04835_),
    .Z(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10129_ (.I(_04838_),
    .Z(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10130_ (.I0(_04817_),
    .I1(\u2.mem[46][15] ),
    .S(_04835_),
    .Z(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10131_ (.I(_04839_),
    .Z(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10132_ (.A1(_04417_),
    .A2(_04760_),
    .ZN(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10133_ (.I(_04840_),
    .Z(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10134_ (.I0(_04782_),
    .I1(\u2.mem[47][0] ),
    .S(_04841_),
    .Z(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10135_ (.I(_04842_),
    .Z(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10136_ (.I0(_04786_),
    .I1(\u2.mem[47][1] ),
    .S(_04841_),
    .Z(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10137_ (.I(_04843_),
    .Z(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10138_ (.I0(_04788_),
    .I1(\u2.mem[47][2] ),
    .S(_04841_),
    .Z(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10139_ (.I(_04844_),
    .Z(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10140_ (.I0(_04790_),
    .I1(\u2.mem[47][3] ),
    .S(_04841_),
    .Z(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10141_ (.I(_04845_),
    .Z(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10142_ (.I(_04840_),
    .Z(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10143_ (.I0(_04792_),
    .I1(\u2.mem[47][4] ),
    .S(_04846_),
    .Z(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10144_ (.I(_04847_),
    .Z(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10145_ (.I0(_04795_),
    .I1(\u2.mem[47][5] ),
    .S(_04846_),
    .Z(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10146_ (.I(_04848_),
    .Z(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10147_ (.I0(_04797_),
    .I1(\u2.mem[47][6] ),
    .S(_04846_),
    .Z(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10148_ (.I(_04849_),
    .Z(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10149_ (.I0(_04799_),
    .I1(\u2.mem[47][7] ),
    .S(_04846_),
    .Z(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10150_ (.I(_04850_),
    .Z(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10151_ (.I(_04840_),
    .Z(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10152_ (.I0(_04801_),
    .I1(\u2.mem[47][8] ),
    .S(_04851_),
    .Z(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10153_ (.I(_04852_),
    .Z(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10154_ (.I0(_04804_),
    .I1(\u2.mem[47][9] ),
    .S(_04851_),
    .Z(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10155_ (.I(_04853_),
    .Z(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10156_ (.I0(_04806_),
    .I1(\u2.mem[47][10] ),
    .S(_04851_),
    .Z(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10157_ (.I(_04854_),
    .Z(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10158_ (.I0(_04808_),
    .I1(\u2.mem[47][11] ),
    .S(_04851_),
    .Z(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10159_ (.I(_04855_),
    .Z(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10160_ (.I(_04840_),
    .Z(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10161_ (.I0(_04810_),
    .I1(\u2.mem[47][12] ),
    .S(_04856_),
    .Z(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10162_ (.I(_04857_),
    .Z(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10163_ (.I0(_04813_),
    .I1(\u2.mem[47][13] ),
    .S(_04856_),
    .Z(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10164_ (.I(_04858_),
    .Z(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10165_ (.I0(_04815_),
    .I1(\u2.mem[47][14] ),
    .S(_04856_),
    .Z(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10166_ (.I(_04859_),
    .Z(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10167_ (.I0(_04817_),
    .I1(\u2.mem[47][15] ),
    .S(_04856_),
    .Z(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10168_ (.I(_04860_),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10169_ (.A1(_03477_),
    .A2(\mem_address_trans[5].data_sync ),
    .ZN(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10170_ (.A1(_03478_),
    .A2(_03986_),
    .A3(_04861_),
    .ZN(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10171_ (.I(_04862_),
    .Z(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10172_ (.A1(_03983_),
    .A2(_04863_),
    .ZN(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10173_ (.I(_04864_),
    .Z(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10174_ (.I0(_04782_),
    .I1(\u2.mem[48][0] ),
    .S(_04865_),
    .Z(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10175_ (.I(_04866_),
    .Z(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10176_ (.I0(_04786_),
    .I1(\u2.mem[48][1] ),
    .S(_04865_),
    .Z(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10177_ (.I(_04867_),
    .Z(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10178_ (.I0(_04788_),
    .I1(\u2.mem[48][2] ),
    .S(_04865_),
    .Z(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10179_ (.I(_04868_),
    .Z(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10180_ (.I0(_04790_),
    .I1(\u2.mem[48][3] ),
    .S(_04865_),
    .Z(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10181_ (.I(_04869_),
    .Z(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10182_ (.I(_04864_),
    .Z(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10183_ (.I0(_04792_),
    .I1(\u2.mem[48][4] ),
    .S(_04870_),
    .Z(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10184_ (.I(_04871_),
    .Z(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10185_ (.I0(_04795_),
    .I1(\u2.mem[48][5] ),
    .S(_04870_),
    .Z(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10186_ (.I(_04872_),
    .Z(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10187_ (.I0(_04797_),
    .I1(\u2.mem[48][6] ),
    .S(_04870_),
    .Z(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10188_ (.I(_04873_),
    .Z(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10189_ (.I0(_04799_),
    .I1(\u2.mem[48][7] ),
    .S(_04870_),
    .Z(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10190_ (.I(_04874_),
    .Z(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10191_ (.I(_04864_),
    .Z(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10192_ (.I0(_04801_),
    .I1(\u2.mem[48][8] ),
    .S(_04875_),
    .Z(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10193_ (.I(_04876_),
    .Z(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10194_ (.I0(_04804_),
    .I1(\u2.mem[48][9] ),
    .S(_04875_),
    .Z(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10195_ (.I(_04877_),
    .Z(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10196_ (.I0(_04806_),
    .I1(\u2.mem[48][10] ),
    .S(_04875_),
    .Z(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10197_ (.I(_04878_),
    .Z(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10198_ (.I0(_04808_),
    .I1(\u2.mem[48][11] ),
    .S(_04875_),
    .Z(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10199_ (.I(_04879_),
    .Z(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10200_ (.I(_04864_),
    .Z(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10201_ (.I0(_04810_),
    .I1(\u2.mem[48][12] ),
    .S(_04880_),
    .Z(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10202_ (.I(_04881_),
    .Z(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10203_ (.I0(_04813_),
    .I1(\u2.mem[48][13] ),
    .S(_04880_),
    .Z(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10204_ (.I(_04882_),
    .Z(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10205_ (.I0(_04815_),
    .I1(\u2.mem[48][14] ),
    .S(_04880_),
    .Z(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10206_ (.I(_04883_),
    .Z(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10207_ (.I0(_04817_),
    .I1(\u2.mem[48][15] ),
    .S(_04880_),
    .Z(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10208_ (.I(_04884_),
    .Z(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10209_ (.I(_04564_),
    .Z(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10210_ (.A1(_04013_),
    .A2(_04863_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10211_ (.I(_04886_),
    .Z(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10212_ (.I0(_04885_),
    .I1(\u2.mem[49][0] ),
    .S(_04887_),
    .Z(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10213_ (.I(_04888_),
    .Z(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10214_ (.I(_04569_),
    .Z(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10215_ (.I0(_04889_),
    .I1(\u2.mem[49][1] ),
    .S(_04887_),
    .Z(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10216_ (.I(_04890_),
    .Z(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10217_ (.I(_04572_),
    .Z(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10218_ (.I0(_04891_),
    .I1(\u2.mem[49][2] ),
    .S(_04887_),
    .Z(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10219_ (.I(_04892_),
    .Z(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10220_ (.I(_04575_),
    .Z(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10221_ (.I0(_04893_),
    .I1(\u2.mem[49][3] ),
    .S(_04887_),
    .Z(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10222_ (.I(_04894_),
    .Z(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10223_ (.I(_04578_),
    .Z(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10224_ (.I(_04886_),
    .Z(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10225_ (.I0(_04895_),
    .I1(\u2.mem[49][4] ),
    .S(_04896_),
    .Z(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10226_ (.I(_04897_),
    .Z(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10227_ (.I(_04582_),
    .Z(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10228_ (.I0(_04898_),
    .I1(\u2.mem[49][5] ),
    .S(_04896_),
    .Z(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10229_ (.I(_04899_),
    .Z(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10230_ (.I(_04585_),
    .Z(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10231_ (.I0(_04900_),
    .I1(\u2.mem[49][6] ),
    .S(_04896_),
    .Z(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10232_ (.I(_04901_),
    .Z(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10233_ (.I(_04588_),
    .Z(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10234_ (.I0(_04902_),
    .I1(\u2.mem[49][7] ),
    .S(_04896_),
    .Z(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10235_ (.I(_04903_),
    .Z(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10236_ (.I(_04591_),
    .Z(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10237_ (.I(_04886_),
    .Z(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10238_ (.I0(_04904_),
    .I1(\u2.mem[49][8] ),
    .S(_04905_),
    .Z(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10239_ (.I(_04906_),
    .Z(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10240_ (.I(_04595_),
    .Z(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10241_ (.I0(_04907_),
    .I1(\u2.mem[49][9] ),
    .S(_04905_),
    .Z(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10242_ (.I(_04908_),
    .Z(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10243_ (.I(_04598_),
    .Z(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10244_ (.I0(_04909_),
    .I1(\u2.mem[49][10] ),
    .S(_04905_),
    .Z(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10245_ (.I(_04910_),
    .Z(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10246_ (.I(_04601_),
    .Z(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10247_ (.I0(_04911_),
    .I1(\u2.mem[49][11] ),
    .S(_04905_),
    .Z(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10248_ (.I(_04912_),
    .Z(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10249_ (.I(_04604_),
    .Z(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10250_ (.I(_04886_),
    .Z(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10251_ (.I0(_04913_),
    .I1(\u2.mem[49][12] ),
    .S(_04914_),
    .Z(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10252_ (.I(_04915_),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10253_ (.I(_04608_),
    .Z(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10254_ (.I0(_04916_),
    .I1(\u2.mem[49][13] ),
    .S(_04914_),
    .Z(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10255_ (.I(_04917_),
    .Z(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10256_ (.I(_04611_),
    .Z(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10257_ (.I0(_04918_),
    .I1(\u2.mem[49][14] ),
    .S(_04914_),
    .Z(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10258_ (.I(_04919_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10259_ (.I(_04614_),
    .Z(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10260_ (.I0(_04920_),
    .I1(\u2.mem[49][15] ),
    .S(_04914_),
    .Z(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10261_ (.I(_04921_),
    .Z(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10262_ (.A1(_03583_),
    .A2(_04863_),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10263_ (.I(_04922_),
    .Z(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10264_ (.I0(_04885_),
    .I1(\u2.mem[50][0] ),
    .S(_04923_),
    .Z(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10265_ (.I(_04924_),
    .Z(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10266_ (.I0(_04889_),
    .I1(\u2.mem[50][1] ),
    .S(_04923_),
    .Z(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10267_ (.I(_04925_),
    .Z(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10268_ (.I0(_04891_),
    .I1(\u2.mem[50][2] ),
    .S(_04923_),
    .Z(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10269_ (.I(_04926_),
    .Z(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10270_ (.I0(_04893_),
    .I1(\u2.mem[50][3] ),
    .S(_04923_),
    .Z(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10271_ (.I(_04927_),
    .Z(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10272_ (.I(_04922_),
    .Z(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10273_ (.I0(_04895_),
    .I1(\u2.mem[50][4] ),
    .S(_04928_),
    .Z(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10274_ (.I(_04929_),
    .Z(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10275_ (.I0(_04898_),
    .I1(\u2.mem[50][5] ),
    .S(_04928_),
    .Z(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10276_ (.I(_04930_),
    .Z(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10277_ (.I0(_04900_),
    .I1(\u2.mem[50][6] ),
    .S(_04928_),
    .Z(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10278_ (.I(_04931_),
    .Z(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10279_ (.I0(_04902_),
    .I1(\u2.mem[50][7] ),
    .S(_04928_),
    .Z(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10280_ (.I(_04932_),
    .Z(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10281_ (.I(_04922_),
    .Z(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10282_ (.I0(_04904_),
    .I1(\u2.mem[50][8] ),
    .S(_04933_),
    .Z(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10283_ (.I(_04934_),
    .Z(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10284_ (.I0(_04907_),
    .I1(\u2.mem[50][9] ),
    .S(_04933_),
    .Z(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10285_ (.I(_04935_),
    .Z(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10286_ (.I0(_04909_),
    .I1(\u2.mem[50][10] ),
    .S(_04933_),
    .Z(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10287_ (.I(_04936_),
    .Z(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10288_ (.I0(_04911_),
    .I1(\u2.mem[50][11] ),
    .S(_04933_),
    .Z(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10289_ (.I(_04937_),
    .Z(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10290_ (.I(_04922_),
    .Z(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10291_ (.I0(_04913_),
    .I1(\u2.mem[50][12] ),
    .S(_04938_),
    .Z(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10292_ (.I(_04939_),
    .Z(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10293_ (.I0(_04916_),
    .I1(\u2.mem[50][13] ),
    .S(_04938_),
    .Z(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10294_ (.I(_04940_),
    .Z(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10295_ (.I0(_04918_),
    .I1(\u2.mem[50][14] ),
    .S(_04938_),
    .Z(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10296_ (.I(_04941_),
    .Z(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10297_ (.I0(_04920_),
    .I1(\u2.mem[50][15] ),
    .S(_04938_),
    .Z(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10298_ (.I(_04942_),
    .Z(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10299_ (.A1(_04072_),
    .A2(_04863_),
    .ZN(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10300_ (.I(_04943_),
    .Z(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10301_ (.I0(_04885_),
    .I1(\u2.mem[51][0] ),
    .S(_04944_),
    .Z(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10302_ (.I(_04945_),
    .Z(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10303_ (.I0(_04889_),
    .I1(\u2.mem[51][1] ),
    .S(_04944_),
    .Z(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10304_ (.I(_04946_),
    .Z(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10305_ (.I0(_04891_),
    .I1(\u2.mem[51][2] ),
    .S(_04944_),
    .Z(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10306_ (.I(_04947_),
    .Z(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10307_ (.I0(_04893_),
    .I1(\u2.mem[51][3] ),
    .S(_04944_),
    .Z(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10308_ (.I(_04948_),
    .Z(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10309_ (.I(_04943_),
    .Z(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10310_ (.I0(_04895_),
    .I1(\u2.mem[51][4] ),
    .S(_04949_),
    .Z(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10311_ (.I(_04950_),
    .Z(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10312_ (.I0(_04898_),
    .I1(\u2.mem[51][5] ),
    .S(_04949_),
    .Z(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10313_ (.I(_04951_),
    .Z(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10314_ (.I0(_04900_),
    .I1(\u2.mem[51][6] ),
    .S(_04949_),
    .Z(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10315_ (.I(_04952_),
    .Z(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10316_ (.I0(_04902_),
    .I1(\u2.mem[51][7] ),
    .S(_04949_),
    .Z(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10317_ (.I(_04953_),
    .Z(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10318_ (.I(_04943_),
    .Z(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10319_ (.I0(_04904_),
    .I1(\u2.mem[51][8] ),
    .S(_04954_),
    .Z(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10320_ (.I(_04955_),
    .Z(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10321_ (.I0(_04907_),
    .I1(\u2.mem[51][9] ),
    .S(_04954_),
    .Z(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10322_ (.I(_04956_),
    .Z(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10323_ (.I0(_04909_),
    .I1(\u2.mem[51][10] ),
    .S(_04954_),
    .Z(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10324_ (.I(_04957_),
    .Z(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10325_ (.I0(_04911_),
    .I1(\u2.mem[51][11] ),
    .S(_04954_),
    .Z(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10326_ (.I(_04958_),
    .Z(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10327_ (.I(_04943_),
    .Z(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10328_ (.I0(_04913_),
    .I1(\u2.mem[51][12] ),
    .S(_04959_),
    .Z(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10329_ (.I(_04960_),
    .Z(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10330_ (.I0(_04916_),
    .I1(\u2.mem[51][13] ),
    .S(_04959_),
    .Z(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10331_ (.I(_04961_),
    .Z(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10332_ (.I0(_04918_),
    .I1(\u2.mem[51][14] ),
    .S(_04959_),
    .Z(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10333_ (.I(_04962_),
    .Z(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10334_ (.I0(_04920_),
    .I1(\u2.mem[51][15] ),
    .S(_04959_),
    .Z(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10335_ (.I(_04963_),
    .Z(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10336_ (.I(_04862_),
    .Z(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10337_ (.A1(_04095_),
    .A2(_04964_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10338_ (.I(_04965_),
    .Z(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10339_ (.I0(_04885_),
    .I1(\u2.mem[52][0] ),
    .S(_04966_),
    .Z(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10340_ (.I(_04967_),
    .Z(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10341_ (.I0(_04889_),
    .I1(\u2.mem[52][1] ),
    .S(_04966_),
    .Z(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10342_ (.I(_04968_),
    .Z(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10343_ (.I0(_04891_),
    .I1(\u2.mem[52][2] ),
    .S(_04966_),
    .Z(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10344_ (.I(_04969_),
    .Z(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10345_ (.I0(_04893_),
    .I1(\u2.mem[52][3] ),
    .S(_04966_),
    .Z(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10346_ (.I(_04970_),
    .Z(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10347_ (.I(_04965_),
    .Z(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10348_ (.I0(_04895_),
    .I1(\u2.mem[52][4] ),
    .S(_04971_),
    .Z(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10349_ (.I(_04972_),
    .Z(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10350_ (.I0(_04898_),
    .I1(\u2.mem[52][5] ),
    .S(_04971_),
    .Z(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10351_ (.I(_04973_),
    .Z(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10352_ (.I0(_04900_),
    .I1(\u2.mem[52][6] ),
    .S(_04971_),
    .Z(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10353_ (.I(_04974_),
    .Z(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10354_ (.I0(_04902_),
    .I1(\u2.mem[52][7] ),
    .S(_04971_),
    .Z(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10355_ (.I(_04975_),
    .Z(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10356_ (.I(_04965_),
    .Z(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10357_ (.I0(_04904_),
    .I1(\u2.mem[52][8] ),
    .S(_04976_),
    .Z(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10358_ (.I(_04977_),
    .Z(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10359_ (.I0(_04907_),
    .I1(\u2.mem[52][9] ),
    .S(_04976_),
    .Z(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10360_ (.I(_04978_),
    .Z(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10361_ (.I0(_04909_),
    .I1(\u2.mem[52][10] ),
    .S(_04976_),
    .Z(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10362_ (.I(_04979_),
    .Z(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10363_ (.I0(_04911_),
    .I1(\u2.mem[52][11] ),
    .S(_04976_),
    .Z(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10364_ (.I(_04980_),
    .Z(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10365_ (.I(_04965_),
    .Z(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10366_ (.I0(_04913_),
    .I1(\u2.mem[52][12] ),
    .S(_04981_),
    .Z(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10367_ (.I(_04982_),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10368_ (.I0(_04916_),
    .I1(\u2.mem[52][13] ),
    .S(_04981_),
    .Z(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10369_ (.I(_04983_),
    .Z(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10370_ (.I0(_04918_),
    .I1(\u2.mem[52][14] ),
    .S(_04981_),
    .Z(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10371_ (.I(_04984_),
    .Z(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10372_ (.I0(_04920_),
    .I1(\u2.mem[52][15] ),
    .S(_04981_),
    .Z(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10373_ (.I(_04985_),
    .Z(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10374_ (.I(_04117_),
    .Z(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10375_ (.I(_04986_),
    .Z(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10376_ (.A1(_04121_),
    .A2(_04964_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10377_ (.I(_04988_),
    .Z(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10378_ (.I0(_04987_),
    .I1(\u2.mem[53][0] ),
    .S(_04989_),
    .Z(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10379_ (.I(_04990_),
    .Z(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10380_ (.I(_04126_),
    .Z(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10381_ (.I(_04991_),
    .Z(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10382_ (.I0(_04992_),
    .I1(\u2.mem[53][1] ),
    .S(_04989_),
    .Z(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10383_ (.I(_04993_),
    .Z(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10384_ (.I(_04130_),
    .Z(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10385_ (.I(_04994_),
    .Z(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10386_ (.I0(_04995_),
    .I1(\u2.mem[53][2] ),
    .S(_04989_),
    .Z(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10387_ (.I(_04996_),
    .Z(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10388_ (.I(_04134_),
    .Z(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10389_ (.I(_04997_),
    .Z(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10390_ (.I0(_04998_),
    .I1(\u2.mem[53][3] ),
    .S(_04989_),
    .Z(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10391_ (.I(_04999_),
    .Z(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10392_ (.I(_04138_),
    .Z(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10393_ (.I(_05000_),
    .Z(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10394_ (.I(_04988_),
    .Z(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10395_ (.I0(_05001_),
    .I1(\u2.mem[53][4] ),
    .S(_05002_),
    .Z(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10396_ (.I(_05003_),
    .Z(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10397_ (.I(_04143_),
    .Z(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10398_ (.I(_05004_),
    .Z(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10399_ (.I0(_05005_),
    .I1(\u2.mem[53][5] ),
    .S(_05002_),
    .Z(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10400_ (.I(_05006_),
    .Z(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10401_ (.I(_03683_),
    .Z(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10402_ (.I0(_05007_),
    .I1(\u2.mem[53][6] ),
    .S(_05002_),
    .Z(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10403_ (.I(_05008_),
    .Z(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10404_ (.I(_03687_),
    .Z(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10405_ (.I0(_05009_),
    .I1(\u2.mem[53][7] ),
    .S(_05002_),
    .Z(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10406_ (.I(_05010_),
    .Z(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10407_ (.I(_03691_),
    .Z(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10408_ (.I(_04988_),
    .Z(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10409_ (.I0(_05011_),
    .I1(\u2.mem[53][8] ),
    .S(_05012_),
    .Z(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10410_ (.I(_05013_),
    .Z(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10411_ (.I(_03696_),
    .Z(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10412_ (.I0(_05014_),
    .I1(\u2.mem[53][9] ),
    .S(_05012_),
    .Z(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10413_ (.I(_05015_),
    .Z(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10414_ (.I(_03700_),
    .Z(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10415_ (.I0(_05016_),
    .I1(\u2.mem[53][10] ),
    .S(_05012_),
    .Z(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10416_ (.I(_05017_),
    .Z(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10417_ (.I(_03704_),
    .Z(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10418_ (.I0(_05018_),
    .I1(\u2.mem[53][11] ),
    .S(_05012_),
    .Z(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10419_ (.I(_05019_),
    .Z(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10420_ (.I(_03708_),
    .Z(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10421_ (.I(_04988_),
    .Z(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10422_ (.I0(_05020_),
    .I1(\u2.mem[53][12] ),
    .S(_05021_),
    .Z(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10423_ (.I(_05022_),
    .Z(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10424_ (.I(_03713_),
    .Z(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10425_ (.I0(_05023_),
    .I1(\u2.mem[53][13] ),
    .S(_05021_),
    .Z(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10426_ (.I(_05024_),
    .Z(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10427_ (.I(_03717_),
    .Z(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10428_ (.I0(_05025_),
    .I1(\u2.mem[53][14] ),
    .S(_05021_),
    .Z(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10429_ (.I(_05026_),
    .Z(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10430_ (.I(_03721_),
    .Z(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10431_ (.I0(_05027_),
    .I1(\u2.mem[53][15] ),
    .S(_05021_),
    .Z(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10432_ (.I(_05028_),
    .Z(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10433_ (.A1(_04180_),
    .A2(_04964_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10434_ (.I(_05029_),
    .Z(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10435_ (.I0(_04987_),
    .I1(\u2.mem[54][0] ),
    .S(_05030_),
    .Z(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10436_ (.I(_05031_),
    .Z(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10437_ (.I0(_04992_),
    .I1(\u2.mem[54][1] ),
    .S(_05030_),
    .Z(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10438_ (.I(_05032_),
    .Z(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10439_ (.I0(_04995_),
    .I1(\u2.mem[54][2] ),
    .S(_05030_),
    .Z(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10440_ (.I(_05033_),
    .Z(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10441_ (.I0(_04998_),
    .I1(\u2.mem[54][3] ),
    .S(_05030_),
    .Z(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10442_ (.I(_05034_),
    .Z(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10443_ (.I(_05029_),
    .Z(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10444_ (.I0(_05001_),
    .I1(\u2.mem[54][4] ),
    .S(_05035_),
    .Z(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10445_ (.I(_05036_),
    .Z(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10446_ (.I0(_05005_),
    .I1(\u2.mem[54][5] ),
    .S(_05035_),
    .Z(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10447_ (.I(_05037_),
    .Z(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10448_ (.I0(_05007_),
    .I1(\u2.mem[54][6] ),
    .S(_05035_),
    .Z(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10449_ (.I(_05038_),
    .Z(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10450_ (.I0(_05009_),
    .I1(\u2.mem[54][7] ),
    .S(_05035_),
    .Z(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10451_ (.I(_05039_),
    .Z(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10452_ (.I(_05029_),
    .Z(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10453_ (.I0(_05011_),
    .I1(\u2.mem[54][8] ),
    .S(_05040_),
    .Z(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10454_ (.I(_05041_),
    .Z(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10455_ (.I0(_05014_),
    .I1(\u2.mem[54][9] ),
    .S(_05040_),
    .Z(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10456_ (.I(_05042_),
    .Z(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10457_ (.I0(_05016_),
    .I1(\u2.mem[54][10] ),
    .S(_05040_),
    .Z(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10458_ (.I(_05043_),
    .Z(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10459_ (.I0(_05018_),
    .I1(\u2.mem[54][11] ),
    .S(_05040_),
    .Z(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10460_ (.I(_05044_),
    .Z(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10461_ (.I(_05029_),
    .Z(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10462_ (.I0(_05020_),
    .I1(\u2.mem[54][12] ),
    .S(_05045_),
    .Z(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10463_ (.I(_05046_),
    .Z(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10464_ (.I0(_05023_),
    .I1(\u2.mem[54][13] ),
    .S(_05045_),
    .Z(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10465_ (.I(_05047_),
    .Z(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10466_ (.I0(_05025_),
    .I1(\u2.mem[54][14] ),
    .S(_05045_),
    .Z(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10467_ (.I(_05048_),
    .Z(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10468_ (.I0(_05027_),
    .I1(\u2.mem[54][15] ),
    .S(_05045_),
    .Z(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10469_ (.I(_05049_),
    .Z(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10470_ (.A1(_03752_),
    .A2(_04964_),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10471_ (.I(_05050_),
    .Z(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10472_ (.I0(_04987_),
    .I1(\u2.mem[55][0] ),
    .S(_05051_),
    .Z(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10473_ (.I(_05052_),
    .Z(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10474_ (.I0(_04992_),
    .I1(\u2.mem[55][1] ),
    .S(_05051_),
    .Z(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10475_ (.I(_05053_),
    .Z(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10476_ (.I0(_04995_),
    .I1(\u2.mem[55][2] ),
    .S(_05051_),
    .Z(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10477_ (.I(_05054_),
    .Z(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10478_ (.I0(_04998_),
    .I1(\u2.mem[55][3] ),
    .S(_05051_),
    .Z(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10479_ (.I(_05055_),
    .Z(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10480_ (.I(_05050_),
    .Z(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10481_ (.I0(_05001_),
    .I1(\u2.mem[55][4] ),
    .S(_05056_),
    .Z(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10482_ (.I(_05057_),
    .Z(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10483_ (.I0(_05005_),
    .I1(\u2.mem[55][5] ),
    .S(_05056_),
    .Z(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10484_ (.I(_05058_),
    .Z(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10485_ (.I0(_05007_),
    .I1(\u2.mem[55][6] ),
    .S(_05056_),
    .Z(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10486_ (.I(_05059_),
    .Z(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10487_ (.I0(_05009_),
    .I1(\u2.mem[55][7] ),
    .S(_05056_),
    .Z(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10488_ (.I(_05060_),
    .Z(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10489_ (.I(_05050_),
    .Z(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10490_ (.I0(_05011_),
    .I1(\u2.mem[55][8] ),
    .S(_05061_),
    .Z(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10491_ (.I(_05062_),
    .Z(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10492_ (.I0(_05014_),
    .I1(\u2.mem[55][9] ),
    .S(_05061_),
    .Z(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10493_ (.I(_05063_),
    .Z(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10494_ (.I0(_05016_),
    .I1(\u2.mem[55][10] ),
    .S(_05061_),
    .Z(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10495_ (.I(_05064_),
    .Z(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10496_ (.I0(_05018_),
    .I1(\u2.mem[55][11] ),
    .S(_05061_),
    .Z(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10497_ (.I(_05065_),
    .Z(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10498_ (.I(_05050_),
    .Z(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10499_ (.I0(_05020_),
    .I1(\u2.mem[55][12] ),
    .S(_05066_),
    .Z(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10500_ (.I(_05067_),
    .Z(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10501_ (.I0(_05023_),
    .I1(\u2.mem[55][13] ),
    .S(_05066_),
    .Z(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10502_ (.I(_05068_),
    .Z(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10503_ (.I0(_05025_),
    .I1(\u2.mem[55][14] ),
    .S(_05066_),
    .Z(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10504_ (.I(_05069_),
    .Z(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10505_ (.I0(_05027_),
    .I1(\u2.mem[55][15] ),
    .S(_05066_),
    .Z(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10506_ (.I(_05070_),
    .Z(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10507_ (.I(_04862_),
    .Z(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10508_ (.A1(_04224_),
    .A2(_05071_),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10509_ (.I(_05072_),
    .Z(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10510_ (.I0(_04987_),
    .I1(\u2.mem[56][0] ),
    .S(_05073_),
    .Z(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10511_ (.I(_05074_),
    .Z(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10512_ (.I0(_04992_),
    .I1(\u2.mem[56][1] ),
    .S(_05073_),
    .Z(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10513_ (.I(_05075_),
    .Z(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10514_ (.I0(_04995_),
    .I1(\u2.mem[56][2] ),
    .S(_05073_),
    .Z(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10515_ (.I(_05076_),
    .Z(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10516_ (.I0(_04998_),
    .I1(\u2.mem[56][3] ),
    .S(_05073_),
    .Z(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10517_ (.I(_05077_),
    .Z(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10518_ (.I(_05072_),
    .Z(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10519_ (.I0(_05001_),
    .I1(\u2.mem[56][4] ),
    .S(_05078_),
    .Z(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10520_ (.I(_05079_),
    .Z(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10521_ (.I0(_05005_),
    .I1(\u2.mem[56][5] ),
    .S(_05078_),
    .Z(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10522_ (.I(_05080_),
    .Z(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10523_ (.I0(_05007_),
    .I1(\u2.mem[56][6] ),
    .S(_05078_),
    .Z(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10524_ (.I(_05081_),
    .Z(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10525_ (.I0(_05009_),
    .I1(\u2.mem[56][7] ),
    .S(_05078_),
    .Z(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10526_ (.I(_05082_),
    .Z(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10527_ (.I(_05072_),
    .Z(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10528_ (.I0(_05011_),
    .I1(\u2.mem[56][8] ),
    .S(_05083_),
    .Z(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10529_ (.I(_05084_),
    .Z(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10530_ (.I0(_05014_),
    .I1(\u2.mem[56][9] ),
    .S(_05083_),
    .Z(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10531_ (.I(_05085_),
    .Z(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10532_ (.I0(_05016_),
    .I1(\u2.mem[56][10] ),
    .S(_05083_),
    .Z(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10533_ (.I(_05086_),
    .Z(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10534_ (.I0(_05018_),
    .I1(\u2.mem[56][11] ),
    .S(_05083_),
    .Z(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10535_ (.I(_05087_),
    .Z(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10536_ (.I(_05072_),
    .Z(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10537_ (.I0(_05020_),
    .I1(\u2.mem[56][12] ),
    .S(_05088_),
    .Z(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10538_ (.I(_05089_),
    .Z(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10539_ (.I0(_05023_),
    .I1(\u2.mem[56][13] ),
    .S(_05088_),
    .Z(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10540_ (.I(_05090_),
    .Z(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10541_ (.I0(_05025_),
    .I1(\u2.mem[56][14] ),
    .S(_05088_),
    .Z(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10542_ (.I(_05091_),
    .Z(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10543_ (.I0(_05027_),
    .I1(\u2.mem[56][15] ),
    .S(_05088_),
    .Z(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10544_ (.I(_05092_),
    .Z(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10545_ (.I(_04986_),
    .Z(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10546_ (.A1(_04249_),
    .A2(_05071_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10547_ (.I(_05094_),
    .Z(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10548_ (.I0(_05093_),
    .I1(\u2.mem[57][0] ),
    .S(_05095_),
    .Z(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10549_ (.I(_05096_),
    .Z(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10550_ (.I(_04991_),
    .Z(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10551_ (.I0(_05097_),
    .I1(\u2.mem[57][1] ),
    .S(_05095_),
    .Z(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10552_ (.I(_05098_),
    .Z(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10553_ (.I(_04994_),
    .Z(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10554_ (.I0(_05099_),
    .I1(\u2.mem[57][2] ),
    .S(_05095_),
    .Z(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10555_ (.I(_05100_),
    .Z(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10556_ (.I(_04997_),
    .Z(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10557_ (.I0(_05101_),
    .I1(\u2.mem[57][3] ),
    .S(_05095_),
    .Z(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10558_ (.I(_05102_),
    .Z(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10559_ (.I(_05000_),
    .Z(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10560_ (.I(_05094_),
    .Z(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10561_ (.I0(_05103_),
    .I1(\u2.mem[57][4] ),
    .S(_05104_),
    .Z(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10562_ (.I(_05105_),
    .Z(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10563_ (.I(_05004_),
    .Z(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10564_ (.I0(_05106_),
    .I1(\u2.mem[57][5] ),
    .S(_05104_),
    .Z(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10565_ (.I(_05107_),
    .Z(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10566_ (.I(_03683_),
    .Z(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10567_ (.I0(_05108_),
    .I1(\u2.mem[57][6] ),
    .S(_05104_),
    .Z(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10568_ (.I(_05109_),
    .Z(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10569_ (.I(_03687_),
    .Z(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10570_ (.I0(_05110_),
    .I1(\u2.mem[57][7] ),
    .S(_05104_),
    .Z(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10571_ (.I(_05111_),
    .Z(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10572_ (.I(_03691_),
    .Z(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10573_ (.I(_05094_),
    .Z(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10574_ (.I0(_05112_),
    .I1(\u2.mem[57][8] ),
    .S(_05113_),
    .Z(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10575_ (.I(_05114_),
    .Z(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10576_ (.I(_03696_),
    .Z(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10577_ (.I0(_05115_),
    .I1(\u2.mem[57][9] ),
    .S(_05113_),
    .Z(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10578_ (.I(_05116_),
    .Z(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10579_ (.I(_03700_),
    .Z(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10580_ (.I0(_05117_),
    .I1(\u2.mem[57][10] ),
    .S(_05113_),
    .Z(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10581_ (.I(_05118_),
    .Z(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10582_ (.I(_03704_),
    .Z(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10583_ (.I0(_05119_),
    .I1(\u2.mem[57][11] ),
    .S(_05113_),
    .Z(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10584_ (.I(_05120_),
    .Z(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10585_ (.I(_03708_),
    .Z(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10586_ (.I(_05094_),
    .Z(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10587_ (.I0(_05121_),
    .I1(\u2.mem[57][12] ),
    .S(_05122_),
    .Z(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10588_ (.I(_05123_),
    .Z(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10589_ (.I(_03713_),
    .Z(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10590_ (.I0(_05124_),
    .I1(\u2.mem[57][13] ),
    .S(_05122_),
    .Z(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10591_ (.I(_05125_),
    .Z(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10592_ (.I(_03717_),
    .Z(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10593_ (.I0(_05126_),
    .I1(\u2.mem[57][14] ),
    .S(_05122_),
    .Z(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10594_ (.I(_05127_),
    .Z(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10595_ (.I(_03721_),
    .Z(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10596_ (.I0(_05128_),
    .I1(\u2.mem[57][15] ),
    .S(_05122_),
    .Z(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10597_ (.I(_05129_),
    .Z(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10598_ (.A1(_04288_),
    .A2(_05071_),
    .ZN(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10599_ (.I(_05130_),
    .Z(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10600_ (.I0(_05093_),
    .I1(\u2.mem[58][0] ),
    .S(_05131_),
    .Z(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10601_ (.I(_05132_),
    .Z(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10602_ (.I0(_05097_),
    .I1(\u2.mem[58][1] ),
    .S(_05131_),
    .Z(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10603_ (.I(_05133_),
    .Z(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10604_ (.I0(_05099_),
    .I1(\u2.mem[58][2] ),
    .S(_05131_),
    .Z(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10605_ (.I(_05134_),
    .Z(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10606_ (.I0(_05101_),
    .I1(\u2.mem[58][3] ),
    .S(_05131_),
    .Z(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10607_ (.I(_05135_),
    .Z(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10608_ (.I(_05130_),
    .Z(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10609_ (.I0(_05103_),
    .I1(\u2.mem[58][4] ),
    .S(_05136_),
    .Z(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10610_ (.I(_05137_),
    .Z(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10611_ (.I0(_05106_),
    .I1(\u2.mem[58][5] ),
    .S(_05136_),
    .Z(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10612_ (.I(_05138_),
    .Z(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10613_ (.I0(_05108_),
    .I1(\u2.mem[58][6] ),
    .S(_05136_),
    .Z(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10614_ (.I(_05139_),
    .Z(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10615_ (.I0(_05110_),
    .I1(\u2.mem[58][7] ),
    .S(_05136_),
    .Z(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10616_ (.I(_05140_),
    .Z(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10617_ (.I(_05130_),
    .Z(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10618_ (.I0(_05112_),
    .I1(\u2.mem[58][8] ),
    .S(_05141_),
    .Z(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10619_ (.I(_05142_),
    .Z(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10620_ (.I0(_05115_),
    .I1(\u2.mem[58][9] ),
    .S(_05141_),
    .Z(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10621_ (.I(_05143_),
    .Z(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10622_ (.I0(_05117_),
    .I1(\u2.mem[58][10] ),
    .S(_05141_),
    .Z(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10623_ (.I(_05144_),
    .Z(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10624_ (.I0(_05119_),
    .I1(\u2.mem[58][11] ),
    .S(_05141_),
    .Z(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10625_ (.I(_05145_),
    .Z(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10626_ (.I(_05130_),
    .Z(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10627_ (.I0(_05121_),
    .I1(\u2.mem[58][12] ),
    .S(_05146_),
    .Z(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10628_ (.I(_05147_),
    .Z(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10629_ (.I0(_05124_),
    .I1(\u2.mem[58][13] ),
    .S(_05146_),
    .Z(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10630_ (.I(_05148_),
    .Z(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10631_ (.I0(_05126_),
    .I1(\u2.mem[58][14] ),
    .S(_05146_),
    .Z(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10632_ (.I(_05149_),
    .Z(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10633_ (.I0(_05128_),
    .I1(\u2.mem[58][15] ),
    .S(_05146_),
    .Z(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10634_ (.I(_05150_),
    .Z(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10635_ (.A1(_04311_),
    .A2(_05071_),
    .ZN(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10636_ (.I(_05151_),
    .Z(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10637_ (.I0(_05093_),
    .I1(\u2.mem[59][0] ),
    .S(_05152_),
    .Z(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10638_ (.I(_05153_),
    .Z(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10639_ (.I0(_05097_),
    .I1(\u2.mem[59][1] ),
    .S(_05152_),
    .Z(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10640_ (.I(_05154_),
    .Z(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10641_ (.I0(_05099_),
    .I1(\u2.mem[59][2] ),
    .S(_05152_),
    .Z(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10642_ (.I(_05155_),
    .Z(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10643_ (.I0(_05101_),
    .I1(\u2.mem[59][3] ),
    .S(_05152_),
    .Z(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10644_ (.I(_05156_),
    .Z(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10645_ (.I(_05151_),
    .Z(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10646_ (.I0(_05103_),
    .I1(\u2.mem[59][4] ),
    .S(_05157_),
    .Z(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10647_ (.I(_05158_),
    .Z(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10648_ (.I0(_05106_),
    .I1(\u2.mem[59][5] ),
    .S(_05157_),
    .Z(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10649_ (.I(_05159_),
    .Z(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10650_ (.I0(_05108_),
    .I1(\u2.mem[59][6] ),
    .S(_05157_),
    .Z(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10651_ (.I(_05160_),
    .Z(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10652_ (.I0(_05110_),
    .I1(\u2.mem[59][7] ),
    .S(_05157_),
    .Z(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10653_ (.I(_05161_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10654_ (.I(_05151_),
    .Z(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10655_ (.I0(_05112_),
    .I1(\u2.mem[59][8] ),
    .S(_05162_),
    .Z(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10656_ (.I(_05163_),
    .Z(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10657_ (.I0(_05115_),
    .I1(\u2.mem[59][9] ),
    .S(_05162_),
    .Z(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10658_ (.I(_05164_),
    .Z(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10659_ (.I0(_05117_),
    .I1(\u2.mem[59][10] ),
    .S(_05162_),
    .Z(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10660_ (.I(_05165_),
    .Z(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10661_ (.I0(_05119_),
    .I1(\u2.mem[59][11] ),
    .S(_05162_),
    .Z(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10662_ (.I(_05166_),
    .Z(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10663_ (.I(_05151_),
    .Z(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10664_ (.I0(_05121_),
    .I1(\u2.mem[59][12] ),
    .S(_05167_),
    .Z(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10665_ (.I(_05168_),
    .Z(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10666_ (.I0(_05124_),
    .I1(\u2.mem[59][13] ),
    .S(_05167_),
    .Z(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10667_ (.I(_05169_),
    .Z(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10668_ (.I0(_05126_),
    .I1(\u2.mem[59][14] ),
    .S(_05167_),
    .Z(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10669_ (.I(_05170_),
    .Z(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10670_ (.I0(_05128_),
    .I1(\u2.mem[59][15] ),
    .S(_05167_),
    .Z(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10671_ (.I(_05171_),
    .Z(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10672_ (.I(_04862_),
    .Z(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10673_ (.A1(_04334_),
    .A2(_05172_),
    .ZN(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10674_ (.I(_05173_),
    .Z(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10675_ (.I0(_05093_),
    .I1(\u2.mem[60][0] ),
    .S(_05174_),
    .Z(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10676_ (.I(_05175_),
    .Z(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10677_ (.I0(_05097_),
    .I1(\u2.mem[60][1] ),
    .S(_05174_),
    .Z(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10678_ (.I(_05176_),
    .Z(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10679_ (.I0(_05099_),
    .I1(\u2.mem[60][2] ),
    .S(_05174_),
    .Z(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10680_ (.I(_05177_),
    .Z(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10681_ (.I0(_05101_),
    .I1(\u2.mem[60][3] ),
    .S(_05174_),
    .Z(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10682_ (.I(_05178_),
    .Z(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10683_ (.I(_05173_),
    .Z(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10684_ (.I0(_05103_),
    .I1(\u2.mem[60][4] ),
    .S(_05179_),
    .Z(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10685_ (.I(_05180_),
    .Z(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10686_ (.I0(_05106_),
    .I1(\u2.mem[60][5] ),
    .S(_05179_),
    .Z(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10687_ (.I(_05181_),
    .Z(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10688_ (.I0(_05108_),
    .I1(\u2.mem[60][6] ),
    .S(_05179_),
    .Z(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10689_ (.I(_05182_),
    .Z(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10690_ (.I0(_05110_),
    .I1(\u2.mem[60][7] ),
    .S(_05179_),
    .Z(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10691_ (.I(_05183_),
    .Z(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10692_ (.I(_05173_),
    .Z(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10693_ (.I0(_05112_),
    .I1(\u2.mem[60][8] ),
    .S(_05184_),
    .Z(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10694_ (.I(_05185_),
    .Z(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10695_ (.I0(_05115_),
    .I1(\u2.mem[60][9] ),
    .S(_05184_),
    .Z(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10696_ (.I(_05186_),
    .Z(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10697_ (.I0(_05117_),
    .I1(\u2.mem[60][10] ),
    .S(_05184_),
    .Z(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10698_ (.I(_05187_),
    .Z(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10699_ (.I0(_05119_),
    .I1(\u2.mem[60][11] ),
    .S(_05184_),
    .Z(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10700_ (.I(_05188_),
    .Z(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10701_ (.I(_05173_),
    .Z(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10702_ (.I0(_05121_),
    .I1(\u2.mem[60][12] ),
    .S(_05189_),
    .Z(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10703_ (.I(_05190_),
    .Z(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10704_ (.I0(_05124_),
    .I1(\u2.mem[60][13] ),
    .S(_05189_),
    .Z(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10705_ (.I(_05191_),
    .Z(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10706_ (.I0(_05126_),
    .I1(\u2.mem[60][14] ),
    .S(_05189_),
    .Z(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10707_ (.I(_05192_),
    .Z(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10708_ (.I0(_05128_),
    .I1(\u2.mem[60][15] ),
    .S(_05189_),
    .Z(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10709_ (.I(_05193_),
    .Z(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10710_ (.I(_04986_),
    .Z(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10711_ (.A1(_03904_),
    .A2(_05172_),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10712_ (.I(_05195_),
    .Z(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10713_ (.I0(_05194_),
    .I1(\u2.mem[61][0] ),
    .S(_05196_),
    .Z(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10714_ (.I(_05197_),
    .Z(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10715_ (.I(_04991_),
    .Z(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10716_ (.I0(_05198_),
    .I1(\u2.mem[61][1] ),
    .S(_05196_),
    .Z(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10717_ (.I(_05199_),
    .Z(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10718_ (.I(_04994_),
    .Z(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10719_ (.I0(_05200_),
    .I1(\u2.mem[61][2] ),
    .S(_05196_),
    .Z(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10720_ (.I(_05201_),
    .Z(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10721_ (.I(_04997_),
    .Z(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10722_ (.I0(_05202_),
    .I1(\u2.mem[61][3] ),
    .S(_05196_),
    .Z(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10723_ (.I(_05203_),
    .Z(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10724_ (.I(_05000_),
    .Z(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10725_ (.I(_05195_),
    .Z(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10726_ (.I0(_05204_),
    .I1(\u2.mem[61][4] ),
    .S(_05205_),
    .Z(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10727_ (.I(_05206_),
    .Z(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10728_ (.I(_05004_),
    .Z(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10729_ (.I0(_05207_),
    .I1(\u2.mem[61][5] ),
    .S(_05205_),
    .Z(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10730_ (.I(_05208_),
    .Z(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10731_ (.I(_03683_),
    .Z(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10732_ (.I0(_05209_),
    .I1(\u2.mem[61][6] ),
    .S(_05205_),
    .Z(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10733_ (.I(_05210_),
    .Z(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10734_ (.I(_03687_),
    .Z(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10735_ (.I0(_05211_),
    .I1(\u2.mem[61][7] ),
    .S(_05205_),
    .Z(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10736_ (.I(_05212_),
    .Z(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10737_ (.I(_03691_),
    .Z(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10738_ (.I(_05195_),
    .Z(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10739_ (.I0(_05213_),
    .I1(\u2.mem[61][8] ),
    .S(_05214_),
    .Z(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10740_ (.I(_05215_),
    .Z(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10741_ (.I(_03696_),
    .Z(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10742_ (.I0(_05216_),
    .I1(\u2.mem[61][9] ),
    .S(_05214_),
    .Z(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10743_ (.I(_05217_),
    .Z(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10744_ (.I(_03700_),
    .Z(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10745_ (.I0(_05218_),
    .I1(\u2.mem[61][10] ),
    .S(_05214_),
    .Z(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10746_ (.I(_05219_),
    .Z(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10747_ (.I(_03704_),
    .Z(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10748_ (.I0(_05220_),
    .I1(\u2.mem[61][11] ),
    .S(_05214_),
    .Z(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10749_ (.I(_05221_),
    .Z(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10750_ (.I(_03708_),
    .Z(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10751_ (.I(_05195_),
    .Z(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10752_ (.I0(_05222_),
    .I1(\u2.mem[61][12] ),
    .S(_05223_),
    .Z(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10753_ (.I(_05224_),
    .Z(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10754_ (.I(_03713_),
    .Z(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10755_ (.I0(_05225_),
    .I1(\u2.mem[61][13] ),
    .S(_05223_),
    .Z(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10756_ (.I(_05226_),
    .Z(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10757_ (.I(_03717_),
    .Z(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10758_ (.I0(_05227_),
    .I1(\u2.mem[61][14] ),
    .S(_05223_),
    .Z(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10759_ (.I(_05228_),
    .Z(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10760_ (.I(_03721_),
    .Z(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10761_ (.I0(_05229_),
    .I1(\u2.mem[61][15] ),
    .S(_05223_),
    .Z(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10762_ (.I(_05230_),
    .Z(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10763_ (.A1(_04394_),
    .A2(_05172_),
    .ZN(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10764_ (.I(_05231_),
    .Z(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10765_ (.I0(_05194_),
    .I1(\u2.mem[62][0] ),
    .S(_05232_),
    .Z(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10766_ (.I(_05233_),
    .Z(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10767_ (.I0(_05198_),
    .I1(\u2.mem[62][1] ),
    .S(_05232_),
    .Z(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10768_ (.I(_05234_),
    .Z(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10769_ (.I0(_05200_),
    .I1(\u2.mem[62][2] ),
    .S(_05232_),
    .Z(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10770_ (.I(_05235_),
    .Z(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10771_ (.I0(_05202_),
    .I1(\u2.mem[62][3] ),
    .S(_05232_),
    .Z(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10772_ (.I(_05236_),
    .Z(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10773_ (.I(_05231_),
    .Z(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10774_ (.I0(_05204_),
    .I1(\u2.mem[62][4] ),
    .S(_05237_),
    .Z(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10775_ (.I(_05238_),
    .Z(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10776_ (.I0(_05207_),
    .I1(\u2.mem[62][5] ),
    .S(_05237_),
    .Z(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10777_ (.I(_05239_),
    .Z(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10778_ (.I0(_05209_),
    .I1(\u2.mem[62][6] ),
    .S(_05237_),
    .Z(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10779_ (.I(_05240_),
    .Z(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10780_ (.I0(_05211_),
    .I1(\u2.mem[62][7] ),
    .S(_05237_),
    .Z(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10781_ (.I(_05241_),
    .Z(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10782_ (.I(_05231_),
    .Z(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10783_ (.I0(_05213_),
    .I1(\u2.mem[62][8] ),
    .S(_05242_),
    .Z(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10784_ (.I(_05243_),
    .Z(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10785_ (.I0(_05216_),
    .I1(\u2.mem[62][9] ),
    .S(_05242_),
    .Z(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10786_ (.I(_05244_),
    .Z(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10787_ (.I0(_05218_),
    .I1(\u2.mem[62][10] ),
    .S(_05242_),
    .Z(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10788_ (.I(_05245_),
    .Z(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10789_ (.I0(_05220_),
    .I1(\u2.mem[62][11] ),
    .S(_05242_),
    .Z(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10790_ (.I(_05246_),
    .Z(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10791_ (.I(_05231_),
    .Z(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10792_ (.I0(_05222_),
    .I1(\u2.mem[62][12] ),
    .S(_05247_),
    .Z(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10793_ (.I(_05248_),
    .Z(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10794_ (.I0(_05225_),
    .I1(\u2.mem[62][13] ),
    .S(_05247_),
    .Z(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10795_ (.I(_05249_),
    .Z(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10796_ (.I0(_05227_),
    .I1(\u2.mem[62][14] ),
    .S(_05247_),
    .Z(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10797_ (.I(_05250_),
    .Z(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10798_ (.I0(_05229_),
    .I1(\u2.mem[62][15] ),
    .S(_05247_),
    .Z(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10799_ (.I(_05251_),
    .Z(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10800_ (.A1(_04416_),
    .A2(_05172_),
    .Z(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10801_ (.I(_05252_),
    .Z(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10802_ (.I0(\u2.mem[63][0] ),
    .I1(_03492_),
    .S(_05253_),
    .Z(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10803_ (.I(_05254_),
    .Z(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10804_ (.I0(\u2.mem[63][1] ),
    .I1(_03497_),
    .S(_05253_),
    .Z(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10805_ (.I(_05255_),
    .Z(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10806_ (.I0(\u2.mem[63][2] ),
    .I1(_03500_),
    .S(_05253_),
    .Z(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10807_ (.I(_05256_),
    .Z(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10808_ (.I0(\u2.mem[63][3] ),
    .I1(_03503_),
    .S(_05253_),
    .Z(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10809_ (.I(_05257_),
    .Z(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10810_ (.I(_05252_),
    .Z(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10811_ (.I0(\u2.mem[63][4] ),
    .I1(_03507_),
    .S(_05258_),
    .Z(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10812_ (.I(_05259_),
    .Z(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10813_ (.I0(\u2.mem[63][5] ),
    .I1(_03511_),
    .S(_05258_),
    .Z(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10814_ (.I(_05260_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10815_ (.I0(\u2.mem[63][6] ),
    .I1(_03513_),
    .S(_05258_),
    .Z(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10816_ (.I(_05261_),
    .Z(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10817_ (.I0(\u2.mem[63][7] ),
    .I1(_03515_),
    .S(_05258_),
    .Z(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10818_ (.I(_05262_),
    .Z(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10819_ (.I(_05252_),
    .Z(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10820_ (.I0(\u2.mem[63][8] ),
    .I1(_03518_),
    .S(_05263_),
    .Z(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10821_ (.I(_05264_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10822_ (.I0(\u2.mem[63][9] ),
    .I1(_03521_),
    .S(_05263_),
    .Z(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10823_ (.I(_05265_),
    .Z(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10824_ (.I0(\u2.mem[63][10] ),
    .I1(_03523_),
    .S(_05263_),
    .Z(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10825_ (.I(_05266_),
    .Z(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10826_ (.I0(\u2.mem[63][11] ),
    .I1(_03525_),
    .S(_05263_),
    .Z(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10827_ (.I(_05267_),
    .Z(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10828_ (.I(_05252_),
    .Z(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10829_ (.I0(\u2.mem[63][12] ),
    .I1(_03528_),
    .S(_05268_),
    .Z(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10830_ (.I(_05269_),
    .Z(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10831_ (.I0(\u2.mem[63][13] ),
    .I1(_03531_),
    .S(_05268_),
    .Z(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10832_ (.I(_05270_),
    .Z(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10833_ (.I0(\u2.mem[63][14] ),
    .I1(_03533_),
    .S(_05268_),
    .Z(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10834_ (.I(_05271_),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10835_ (.I0(\u2.mem[63][15] ),
    .I1(_05229_),
    .S(_05268_),
    .Z(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10836_ (.I(_05272_),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10837_ (.I(\mem_address_trans[6].data_sync ),
    .ZN(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10838_ (.A1(_05273_),
    .A2(_03986_),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10839_ (.A1(_03477_),
    .A2(_03985_),
    .A3(_05274_),
    .ZN(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10840_ (.I(_05275_),
    .Z(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10841_ (.A1(_03983_),
    .A2(_05276_),
    .ZN(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10842_ (.I(_05277_),
    .Z(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10843_ (.I0(_05194_),
    .I1(\u2.mem[128][0] ),
    .S(_05278_),
    .Z(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10844_ (.I(_05279_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10845_ (.I0(_05198_),
    .I1(\u2.mem[128][1] ),
    .S(_05278_),
    .Z(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10846_ (.I(_05280_),
    .Z(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10847_ (.I0(_05200_),
    .I1(\u2.mem[128][2] ),
    .S(_05278_),
    .Z(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10848_ (.I(_05281_),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10849_ (.I0(_05202_),
    .I1(\u2.mem[128][3] ),
    .S(_05278_),
    .Z(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10850_ (.I(_05282_),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10851_ (.I0(_05204_),
    .I1(\u2.mem[128][4] ),
    .S(_05277_),
    .Z(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10852_ (.I(_05283_),
    .Z(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10853_ (.I0(_05207_),
    .I1(\u2.mem[128][5] ),
    .S(_05277_),
    .Z(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10854_ (.I(_05284_),
    .Z(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10855_ (.I(_04012_),
    .Z(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10856_ (.A1(_05285_),
    .A2(_05276_),
    .ZN(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10857_ (.I(_05286_),
    .Z(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10858_ (.I0(_05194_),
    .I1(\u2.mem[129][0] ),
    .S(_05287_),
    .Z(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10859_ (.I(_05288_),
    .Z(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10860_ (.I0(_05198_),
    .I1(\u2.mem[129][1] ),
    .S(_05287_),
    .Z(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10861_ (.I(_05289_),
    .Z(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10862_ (.I0(_05200_),
    .I1(\u2.mem[129][2] ),
    .S(_05287_),
    .Z(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10863_ (.I(_05290_),
    .Z(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10864_ (.I0(_05202_),
    .I1(\u2.mem[129][3] ),
    .S(_05287_),
    .Z(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10865_ (.I(_05291_),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10866_ (.I0(_05204_),
    .I1(\u2.mem[129][4] ),
    .S(_05286_),
    .Z(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10867_ (.I(_05292_),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10868_ (.I0(_05207_),
    .I1(\u2.mem[129][5] ),
    .S(_05286_),
    .Z(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10869_ (.I(_05293_),
    .Z(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10870_ (.I(_04986_),
    .Z(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10871_ (.I(_03582_),
    .Z(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10872_ (.A1(_05295_),
    .A2(_05276_),
    .ZN(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10873_ (.I(_05296_),
    .Z(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10874_ (.I0(_05294_),
    .I1(\u2.mem[130][0] ),
    .S(_05297_),
    .Z(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10875_ (.I(_05298_),
    .Z(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10876_ (.I(_04991_),
    .Z(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10877_ (.I0(_05299_),
    .I1(\u2.mem[130][1] ),
    .S(_05297_),
    .Z(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10878_ (.I(_05300_),
    .Z(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10879_ (.I(_04994_),
    .Z(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10880_ (.I0(_05301_),
    .I1(\u2.mem[130][2] ),
    .S(_05297_),
    .Z(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10881_ (.I(_05302_),
    .Z(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10882_ (.I(_04997_),
    .Z(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10883_ (.I0(_05303_),
    .I1(\u2.mem[130][3] ),
    .S(_05297_),
    .Z(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10884_ (.I(_05304_),
    .Z(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10885_ (.I(_05000_),
    .Z(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10886_ (.I0(_05305_),
    .I1(\u2.mem[130][4] ),
    .S(_05296_),
    .Z(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10887_ (.I(_05306_),
    .Z(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10888_ (.I(_05004_),
    .Z(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10889_ (.I0(_05307_),
    .I1(\u2.mem[130][5] ),
    .S(_05296_),
    .Z(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10890_ (.I(_05308_),
    .Z(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10891_ (.A1(_04072_),
    .A2(_05276_),
    .ZN(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10892_ (.I(_05309_),
    .Z(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10893_ (.I0(_05294_),
    .I1(\u2.mem[131][0] ),
    .S(_05310_),
    .Z(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10894_ (.I(_05311_),
    .Z(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10895_ (.I0(_05299_),
    .I1(\u2.mem[131][1] ),
    .S(_05310_),
    .Z(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10896_ (.I(_05312_),
    .Z(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10897_ (.I0(_05301_),
    .I1(\u2.mem[131][2] ),
    .S(_05310_),
    .Z(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10898_ (.I(_05313_),
    .Z(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10899_ (.I0(_05303_),
    .I1(\u2.mem[131][3] ),
    .S(_05310_),
    .Z(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10900_ (.I(_05314_),
    .Z(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10901_ (.I0(_05305_),
    .I1(\u2.mem[131][4] ),
    .S(_05309_),
    .Z(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10902_ (.I(_05315_),
    .Z(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10903_ (.I0(_05307_),
    .I1(\u2.mem[131][5] ),
    .S(_05309_),
    .Z(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10904_ (.I(_05316_),
    .Z(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10905_ (.I(_05275_),
    .Z(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10906_ (.A1(_04095_),
    .A2(_05317_),
    .ZN(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10907_ (.I(_05318_),
    .Z(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10908_ (.I0(_05294_),
    .I1(\u2.mem[132][0] ),
    .S(_05319_),
    .Z(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10909_ (.I(_05320_),
    .Z(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10910_ (.I0(_05299_),
    .I1(\u2.mem[132][1] ),
    .S(_05319_),
    .Z(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10911_ (.I(_05321_),
    .Z(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10912_ (.I0(_05301_),
    .I1(\u2.mem[132][2] ),
    .S(_05319_),
    .Z(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10913_ (.I(_05322_),
    .Z(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10914_ (.I0(_05303_),
    .I1(\u2.mem[132][3] ),
    .S(_05319_),
    .Z(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10915_ (.I(_05323_),
    .Z(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10916_ (.I0(_05305_),
    .I1(\u2.mem[132][4] ),
    .S(_05318_),
    .Z(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10917_ (.I(_05324_),
    .Z(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10918_ (.I0(_05307_),
    .I1(\u2.mem[132][5] ),
    .S(_05318_),
    .Z(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10919_ (.I(_05325_),
    .Z(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10920_ (.A1(_04121_),
    .A2(_05317_),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10921_ (.I(_05326_),
    .Z(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10922_ (.I0(_05294_),
    .I1(\u2.mem[133][0] ),
    .S(_05327_),
    .Z(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10923_ (.I(_05328_),
    .Z(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10924_ (.I0(_05299_),
    .I1(\u2.mem[133][1] ),
    .S(_05327_),
    .Z(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10925_ (.I(_05329_),
    .Z(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10926_ (.I0(_05301_),
    .I1(\u2.mem[133][2] ),
    .S(_05327_),
    .Z(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10927_ (.I(_05330_),
    .Z(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10928_ (.I0(_05303_),
    .I1(\u2.mem[133][3] ),
    .S(_05327_),
    .Z(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10929_ (.I(_05331_),
    .Z(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10930_ (.I0(_05305_),
    .I1(\u2.mem[133][4] ),
    .S(_05326_),
    .Z(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10931_ (.I(_05332_),
    .Z(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10932_ (.I0(_05307_),
    .I1(\u2.mem[133][5] ),
    .S(_05326_),
    .Z(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10933_ (.I(_05333_),
    .Z(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10934_ (.I(_04117_),
    .Z(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10935_ (.I(_05334_),
    .Z(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10936_ (.A1(_04180_),
    .A2(_05317_),
    .ZN(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10937_ (.I(_05336_),
    .Z(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10938_ (.I0(_05335_),
    .I1(\u2.mem[134][0] ),
    .S(_05337_),
    .Z(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10939_ (.I(_05338_),
    .Z(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10940_ (.I(_04126_),
    .Z(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10941_ (.I(_05339_),
    .Z(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10942_ (.I0(_05340_),
    .I1(\u2.mem[134][1] ),
    .S(_05337_),
    .Z(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10943_ (.I(_05341_),
    .Z(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10944_ (.I(_04130_),
    .Z(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10945_ (.I(_05342_),
    .Z(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10946_ (.I0(_05343_),
    .I1(\u2.mem[134][2] ),
    .S(_05337_),
    .Z(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10947_ (.I(_05344_),
    .Z(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10948_ (.I(_04134_),
    .Z(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10949_ (.I(_05345_),
    .Z(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10950_ (.I0(_05346_),
    .I1(\u2.mem[134][3] ),
    .S(_05337_),
    .Z(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10951_ (.I(_05347_),
    .Z(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10952_ (.I(_04138_),
    .Z(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10953_ (.I(_05348_),
    .Z(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10954_ (.I0(_05349_),
    .I1(\u2.mem[134][4] ),
    .S(_05336_),
    .Z(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10955_ (.I(_05350_),
    .Z(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10956_ (.I(_04143_),
    .Z(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10957_ (.I(_05351_),
    .Z(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10958_ (.I0(_05352_),
    .I1(\u2.mem[134][5] ),
    .S(_05336_),
    .Z(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10959_ (.I(_05353_),
    .Z(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10960_ (.I(_03751_),
    .Z(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10961_ (.A1(_05354_),
    .A2(_05317_),
    .ZN(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10962_ (.I(_05355_),
    .Z(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10963_ (.I0(_05335_),
    .I1(\u2.mem[135][0] ),
    .S(_05356_),
    .Z(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10964_ (.I(_05357_),
    .Z(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10965_ (.I0(_05340_),
    .I1(\u2.mem[135][1] ),
    .S(_05356_),
    .Z(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10966_ (.I(_05358_),
    .Z(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10967_ (.I0(_05343_),
    .I1(\u2.mem[135][2] ),
    .S(_05356_),
    .Z(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10968_ (.I(_05359_),
    .Z(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10969_ (.I0(_05346_),
    .I1(\u2.mem[135][3] ),
    .S(_05356_),
    .Z(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10970_ (.I(_05360_),
    .Z(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10971_ (.I0(_05349_),
    .I1(\u2.mem[135][4] ),
    .S(_05355_),
    .Z(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10972_ (.I(_05361_),
    .Z(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10973_ (.I0(_05352_),
    .I1(\u2.mem[135][5] ),
    .S(_05355_),
    .Z(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10974_ (.I(_05362_),
    .Z(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10975_ (.I(_05275_),
    .Z(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10976_ (.A1(_04224_),
    .A2(_05363_),
    .ZN(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10977_ (.I(_05364_),
    .Z(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10978_ (.I0(_05335_),
    .I1(\u2.mem[136][0] ),
    .S(_05365_),
    .Z(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10979_ (.I(_05366_),
    .Z(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10980_ (.I0(_05340_),
    .I1(\u2.mem[136][1] ),
    .S(_05365_),
    .Z(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10981_ (.I(_05367_),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10982_ (.I0(_05343_),
    .I1(\u2.mem[136][2] ),
    .S(_05365_),
    .Z(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10983_ (.I(_05368_),
    .Z(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10984_ (.I0(_05346_),
    .I1(\u2.mem[136][3] ),
    .S(_05365_),
    .Z(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10985_ (.I(_05369_),
    .Z(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10986_ (.I0(_05349_),
    .I1(\u2.mem[136][4] ),
    .S(_05364_),
    .Z(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10987_ (.I(_05370_),
    .Z(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10988_ (.I0(_05352_),
    .I1(\u2.mem[136][5] ),
    .S(_05364_),
    .Z(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10989_ (.I(_05371_),
    .Z(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10990_ (.A1(_04249_),
    .A2(_05363_),
    .ZN(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10991_ (.I(_05372_),
    .Z(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10992_ (.I0(_05335_),
    .I1(\u2.mem[137][0] ),
    .S(_05373_),
    .Z(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10993_ (.I(_05374_),
    .Z(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10994_ (.I0(_05340_),
    .I1(\u2.mem[137][1] ),
    .S(_05373_),
    .Z(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10995_ (.I(_05375_),
    .Z(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10996_ (.I0(_05343_),
    .I1(\u2.mem[137][2] ),
    .S(_05373_),
    .Z(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10997_ (.I(_05376_),
    .Z(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10998_ (.I0(_05346_),
    .I1(\u2.mem[137][3] ),
    .S(_05373_),
    .Z(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10999_ (.I(_05377_),
    .Z(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11000_ (.I0(_05349_),
    .I1(\u2.mem[137][4] ),
    .S(_05372_),
    .Z(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11001_ (.I(_05378_),
    .Z(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11002_ (.I0(_05352_),
    .I1(\u2.mem[137][5] ),
    .S(_05372_),
    .Z(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11003_ (.I(_05379_),
    .Z(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11004_ (.I(_05334_),
    .Z(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11005_ (.A1(_04288_),
    .A2(_05363_),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11006_ (.I(_05381_),
    .Z(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11007_ (.I0(_05380_),
    .I1(\u2.mem[138][0] ),
    .S(_05382_),
    .Z(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11008_ (.I(_05383_),
    .Z(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11009_ (.I(_05339_),
    .Z(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11010_ (.I0(_05384_),
    .I1(\u2.mem[138][1] ),
    .S(_05382_),
    .Z(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11011_ (.I(_05385_),
    .Z(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11012_ (.I(_05342_),
    .Z(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11013_ (.I0(_05386_),
    .I1(\u2.mem[138][2] ),
    .S(_05382_),
    .Z(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11014_ (.I(_05387_),
    .Z(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11015_ (.I(_05345_),
    .Z(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11016_ (.I0(_05388_),
    .I1(\u2.mem[138][3] ),
    .S(_05382_),
    .Z(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11017_ (.I(_05389_),
    .Z(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11018_ (.I(_05348_),
    .Z(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11019_ (.I0(_05390_),
    .I1(\u2.mem[138][4] ),
    .S(_05381_),
    .Z(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11020_ (.I(_05391_),
    .Z(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11021_ (.I(_05351_),
    .Z(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11022_ (.I0(_05392_),
    .I1(\u2.mem[138][5] ),
    .S(_05381_),
    .Z(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11023_ (.I(_05393_),
    .Z(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11024_ (.A1(_04311_),
    .A2(_05363_),
    .ZN(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11025_ (.I(_05394_),
    .Z(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11026_ (.I0(_05380_),
    .I1(\u2.mem[139][0] ),
    .S(_05395_),
    .Z(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11027_ (.I(_05396_),
    .Z(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11028_ (.I0(_05384_),
    .I1(\u2.mem[139][1] ),
    .S(_05395_),
    .Z(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11029_ (.I(_05397_),
    .Z(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11030_ (.I0(_05386_),
    .I1(\u2.mem[139][2] ),
    .S(_05395_),
    .Z(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11031_ (.I(_05398_),
    .Z(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11032_ (.I0(_05388_),
    .I1(\u2.mem[139][3] ),
    .S(_05395_),
    .Z(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11033_ (.I(_05399_),
    .Z(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11034_ (.I0(_05390_),
    .I1(\u2.mem[139][4] ),
    .S(_05394_),
    .Z(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11035_ (.I(_05400_),
    .Z(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11036_ (.I0(_05392_),
    .I1(\u2.mem[139][5] ),
    .S(_05394_),
    .Z(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11037_ (.I(_05401_),
    .Z(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11038_ (.I(_05275_),
    .Z(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11039_ (.A1(_04334_),
    .A2(_05402_),
    .ZN(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11040_ (.I(_05403_),
    .Z(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11041_ (.I0(_05380_),
    .I1(\u2.mem[140][0] ),
    .S(_05404_),
    .Z(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11042_ (.I(_05405_),
    .Z(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11043_ (.I0(_05384_),
    .I1(\u2.mem[140][1] ),
    .S(_05404_),
    .Z(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11044_ (.I(_05406_),
    .Z(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11045_ (.I0(_05386_),
    .I1(\u2.mem[140][2] ),
    .S(_05404_),
    .Z(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11046_ (.I(_05407_),
    .Z(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11047_ (.I0(_05388_),
    .I1(\u2.mem[140][3] ),
    .S(_05404_),
    .Z(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11048_ (.I(_05408_),
    .Z(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11049_ (.I0(_05390_),
    .I1(\u2.mem[140][4] ),
    .S(_05403_),
    .Z(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11050_ (.I(_05409_),
    .Z(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11051_ (.I0(_05392_),
    .I1(\u2.mem[140][5] ),
    .S(_05403_),
    .Z(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11052_ (.I(_05410_),
    .Z(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11053_ (.I(_03903_),
    .Z(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11054_ (.A1(_05411_),
    .A2(_05402_),
    .ZN(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11055_ (.I(_05412_),
    .Z(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11056_ (.I0(_05380_),
    .I1(\u2.mem[141][0] ),
    .S(_05413_),
    .Z(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11057_ (.I(_05414_),
    .Z(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11058_ (.I0(_05384_),
    .I1(\u2.mem[141][1] ),
    .S(_05413_),
    .Z(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11059_ (.I(_05415_),
    .Z(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11060_ (.I0(_05386_),
    .I1(\u2.mem[141][2] ),
    .S(_05413_),
    .Z(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11061_ (.I(_05416_),
    .Z(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11062_ (.I0(_05388_),
    .I1(\u2.mem[141][3] ),
    .S(_05413_),
    .Z(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11063_ (.I(_05417_),
    .Z(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11064_ (.I0(_05390_),
    .I1(\u2.mem[141][4] ),
    .S(_05412_),
    .Z(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11065_ (.I(_05418_),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11066_ (.I0(_05392_),
    .I1(\u2.mem[141][5] ),
    .S(_05412_),
    .Z(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11067_ (.I(_05419_),
    .Z(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11068_ (.I(_05334_),
    .Z(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11069_ (.A1(_04394_),
    .A2(_05402_),
    .ZN(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11070_ (.I(_05421_),
    .Z(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11071_ (.I0(_05420_),
    .I1(\u2.mem[142][0] ),
    .S(_05422_),
    .Z(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11072_ (.I(_05423_),
    .Z(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11073_ (.I(_05339_),
    .Z(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11074_ (.I0(_05424_),
    .I1(\u2.mem[142][1] ),
    .S(_05422_),
    .Z(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11075_ (.I(_05425_),
    .Z(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11076_ (.I(_05342_),
    .Z(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11077_ (.I0(_05426_),
    .I1(\u2.mem[142][2] ),
    .S(_05422_),
    .Z(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11078_ (.I(_05427_),
    .Z(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11079_ (.I(_05345_),
    .Z(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11080_ (.I0(_05428_),
    .I1(\u2.mem[142][3] ),
    .S(_05422_),
    .Z(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11081_ (.I(_05429_),
    .Z(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11082_ (.I(_05348_),
    .Z(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11083_ (.I0(_05430_),
    .I1(\u2.mem[142][4] ),
    .S(_05421_),
    .Z(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11084_ (.I(_05431_),
    .Z(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11085_ (.I(_05351_),
    .Z(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11086_ (.I0(_05432_),
    .I1(\u2.mem[142][5] ),
    .S(_05421_),
    .Z(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11087_ (.I(_05433_),
    .Z(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11088_ (.A1(_04417_),
    .A2(_05402_),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11089_ (.I(_05434_),
    .Z(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11090_ (.I0(_05420_),
    .I1(\u2.mem[143][0] ),
    .S(_05435_),
    .Z(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11091_ (.I(_05436_),
    .Z(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11092_ (.I0(_05424_),
    .I1(\u2.mem[143][1] ),
    .S(_05435_),
    .Z(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11093_ (.I(_05437_),
    .Z(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11094_ (.I0(_05426_),
    .I1(\u2.mem[143][2] ),
    .S(_05435_),
    .Z(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11095_ (.I(_05438_),
    .Z(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11096_ (.I0(_05428_),
    .I1(\u2.mem[143][3] ),
    .S(_05435_),
    .Z(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11097_ (.I(_05439_),
    .Z(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11098_ (.I0(_05430_),
    .I1(\u2.mem[143][4] ),
    .S(_05434_),
    .Z(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11099_ (.I(_05440_),
    .Z(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11100_ (.I0(_05432_),
    .I1(\u2.mem[143][5] ),
    .S(_05434_),
    .Z(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11101_ (.I(_05441_),
    .Z(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _11102_ (.A1(_03984_),
    .A2(_03985_),
    .A3(_05274_),
    .ZN(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11103_ (.I(_05442_),
    .Z(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11104_ (.A1(_03487_),
    .A2(_05443_),
    .ZN(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11105_ (.I(_05444_),
    .Z(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11106_ (.I0(_05420_),
    .I1(\u2.mem[144][0] ),
    .S(_05445_),
    .Z(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11107_ (.I(_05446_),
    .Z(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11108_ (.I0(_05424_),
    .I1(\u2.mem[144][1] ),
    .S(_05445_),
    .Z(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11109_ (.I(_05447_),
    .Z(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11110_ (.I0(_05426_),
    .I1(\u2.mem[144][2] ),
    .S(_05445_),
    .Z(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11111_ (.I(_05448_),
    .Z(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11112_ (.I0(_05428_),
    .I1(\u2.mem[144][3] ),
    .S(_05445_),
    .Z(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11113_ (.I(_05449_),
    .Z(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11114_ (.I0(_05430_),
    .I1(\u2.mem[144][4] ),
    .S(_05444_),
    .Z(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11115_ (.I(_05450_),
    .Z(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11116_ (.I0(_05432_),
    .I1(\u2.mem[144][5] ),
    .S(_05444_),
    .Z(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11117_ (.I(_05451_),
    .Z(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11118_ (.A1(_05285_),
    .A2(_05443_),
    .ZN(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11119_ (.I(_05452_),
    .Z(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11120_ (.I0(_05420_),
    .I1(\u2.mem[145][0] ),
    .S(_05453_),
    .Z(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11121_ (.I(_05454_),
    .Z(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11122_ (.I0(_05424_),
    .I1(\u2.mem[145][1] ),
    .S(_05453_),
    .Z(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11123_ (.I(_05455_),
    .Z(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11124_ (.I0(_05426_),
    .I1(\u2.mem[145][2] ),
    .S(_05453_),
    .Z(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11125_ (.I(_05456_),
    .Z(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11126_ (.I0(_05428_),
    .I1(\u2.mem[145][3] ),
    .S(_05453_),
    .Z(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11127_ (.I(_05457_),
    .Z(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11128_ (.I0(_05430_),
    .I1(\u2.mem[145][4] ),
    .S(_05452_),
    .Z(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11129_ (.I(_05458_),
    .Z(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11130_ (.I0(_05432_),
    .I1(\u2.mem[145][5] ),
    .S(_05452_),
    .Z(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11131_ (.I(_05459_),
    .Z(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11132_ (.I(_05334_),
    .Z(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11133_ (.A1(_05295_),
    .A2(_05443_),
    .ZN(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11134_ (.I(_05461_),
    .Z(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11135_ (.I0(_05460_),
    .I1(\u2.mem[146][0] ),
    .S(_05462_),
    .Z(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11136_ (.I(_05463_),
    .Z(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11137_ (.I(_05339_),
    .Z(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11138_ (.I0(_05464_),
    .I1(\u2.mem[146][1] ),
    .S(_05462_),
    .Z(_05465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11139_ (.I(_05465_),
    .Z(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11140_ (.I(_05342_),
    .Z(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11141_ (.I0(_05466_),
    .I1(\u2.mem[146][2] ),
    .S(_05462_),
    .Z(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11142_ (.I(_05467_),
    .Z(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11143_ (.I(_05345_),
    .Z(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11144_ (.I0(_05468_),
    .I1(\u2.mem[146][3] ),
    .S(_05462_),
    .Z(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11145_ (.I(_05469_),
    .Z(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11146_ (.I(_05348_),
    .Z(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11147_ (.I0(_05470_),
    .I1(\u2.mem[146][4] ),
    .S(_05461_),
    .Z(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11148_ (.I(_05471_),
    .Z(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11149_ (.I(_05351_),
    .Z(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11150_ (.I0(_05472_),
    .I1(\u2.mem[146][5] ),
    .S(_05461_),
    .Z(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11151_ (.I(_05473_),
    .Z(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11152_ (.A1(_04071_),
    .A2(_05443_),
    .ZN(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11153_ (.I(_05474_),
    .Z(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11154_ (.I0(_05460_),
    .I1(\u2.mem[147][0] ),
    .S(_05475_),
    .Z(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11155_ (.I(_05476_),
    .Z(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11156_ (.I0(_05464_),
    .I1(\u2.mem[147][1] ),
    .S(_05475_),
    .Z(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11157_ (.I(_05477_),
    .Z(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11158_ (.I0(_05466_),
    .I1(\u2.mem[147][2] ),
    .S(_05475_),
    .Z(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11159_ (.I(_05478_),
    .Z(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11160_ (.I0(_05468_),
    .I1(\u2.mem[147][3] ),
    .S(_05475_),
    .Z(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11161_ (.I(_05479_),
    .Z(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11162_ (.I0(_05470_),
    .I1(\u2.mem[147][4] ),
    .S(_05474_),
    .Z(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11163_ (.I(_05480_),
    .Z(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11164_ (.I0(_05472_),
    .I1(\u2.mem[147][5] ),
    .S(_05474_),
    .Z(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11165_ (.I(_05481_),
    .Z(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11166_ (.I(_05442_),
    .Z(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11167_ (.A1(_04094_),
    .A2(_05482_),
    .ZN(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11168_ (.I(_05483_),
    .Z(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11169_ (.I0(_05460_),
    .I1(\u2.mem[148][0] ),
    .S(_05484_),
    .Z(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11170_ (.I(_05485_),
    .Z(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11171_ (.I0(_05464_),
    .I1(\u2.mem[148][1] ),
    .S(_05484_),
    .Z(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11172_ (.I(_05486_),
    .Z(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11173_ (.I0(_05466_),
    .I1(\u2.mem[148][2] ),
    .S(_05484_),
    .Z(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11174_ (.I(_05487_),
    .Z(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11175_ (.I0(_05468_),
    .I1(\u2.mem[148][3] ),
    .S(_05484_),
    .Z(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11176_ (.I(_05488_),
    .Z(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11177_ (.I0(_05470_),
    .I1(\u2.mem[148][4] ),
    .S(_05483_),
    .Z(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11178_ (.I(_05489_),
    .Z(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11179_ (.I0(_05472_),
    .I1(\u2.mem[148][5] ),
    .S(_05483_),
    .Z(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11180_ (.I(_05490_),
    .Z(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11181_ (.A1(_04120_),
    .A2(_05482_),
    .ZN(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11182_ (.I(_05491_),
    .Z(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11183_ (.I0(_05460_),
    .I1(\u2.mem[149][0] ),
    .S(_05492_),
    .Z(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11184_ (.I(_05493_),
    .Z(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11185_ (.I0(_05464_),
    .I1(\u2.mem[149][1] ),
    .S(_05492_),
    .Z(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11186_ (.I(_05494_),
    .Z(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11187_ (.I0(_05466_),
    .I1(\u2.mem[149][2] ),
    .S(_05492_),
    .Z(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11188_ (.I(_05495_),
    .Z(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11189_ (.I0(_05468_),
    .I1(\u2.mem[149][3] ),
    .S(_05492_),
    .Z(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11190_ (.I(_05496_),
    .Z(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11191_ (.I0(_05470_),
    .I1(\u2.mem[149][4] ),
    .S(_05491_),
    .Z(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11192_ (.I(_05497_),
    .Z(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11193_ (.I0(_05472_),
    .I1(\u2.mem[149][5] ),
    .S(_05491_),
    .Z(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11194_ (.I(_05498_),
    .Z(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11195_ (.I(_03491_),
    .Z(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11196_ (.I(_05499_),
    .Z(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11197_ (.A1(_04179_),
    .A2(_05482_),
    .ZN(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11198_ (.I(_05501_),
    .Z(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11199_ (.I0(_05500_),
    .I1(\u2.mem[150][0] ),
    .S(_05502_),
    .Z(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11200_ (.I(_05503_),
    .Z(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11201_ (.I(_03496_),
    .Z(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11202_ (.I(_05504_),
    .Z(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11203_ (.I0(_05505_),
    .I1(\u2.mem[150][1] ),
    .S(_05502_),
    .Z(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11204_ (.I(_05506_),
    .Z(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11205_ (.I(_03499_),
    .Z(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11206_ (.I(_05507_),
    .Z(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11207_ (.I0(_05508_),
    .I1(\u2.mem[150][2] ),
    .S(_05502_),
    .Z(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11208_ (.I(_05509_),
    .Z(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11209_ (.I(_03502_),
    .Z(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11210_ (.I(_05510_),
    .Z(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11211_ (.I0(_05511_),
    .I1(\u2.mem[150][3] ),
    .S(_05502_),
    .Z(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11212_ (.I(_05512_),
    .Z(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11213_ (.I(_03506_),
    .Z(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11214_ (.I(_05513_),
    .Z(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11215_ (.I0(_05514_),
    .I1(\u2.mem[150][4] ),
    .S(_05501_),
    .Z(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11216_ (.I(_05515_),
    .Z(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11217_ (.I(_03510_),
    .Z(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11218_ (.I(_05516_),
    .Z(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11219_ (.I0(_05517_),
    .I1(\u2.mem[150][5] ),
    .S(_05501_),
    .Z(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11220_ (.I(_05518_),
    .Z(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11221_ (.A1(_05354_),
    .A2(_05482_),
    .ZN(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11222_ (.I(_05519_),
    .Z(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11223_ (.I0(_05500_),
    .I1(\u2.mem[151][0] ),
    .S(_05520_),
    .Z(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11224_ (.I(_05521_),
    .Z(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11225_ (.I0(_05505_),
    .I1(\u2.mem[151][1] ),
    .S(_05520_),
    .Z(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11226_ (.I(_05522_),
    .Z(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11227_ (.I0(_05508_),
    .I1(\u2.mem[151][2] ),
    .S(_05520_),
    .Z(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11228_ (.I(_05523_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11229_ (.I0(_05511_),
    .I1(\u2.mem[151][3] ),
    .S(_05520_),
    .Z(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11230_ (.I(_05524_),
    .Z(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11231_ (.I0(_05514_),
    .I1(\u2.mem[151][4] ),
    .S(_05519_),
    .Z(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11232_ (.I(_05525_),
    .Z(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11233_ (.I0(_05517_),
    .I1(\u2.mem[151][5] ),
    .S(_05519_),
    .Z(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11234_ (.I(_05526_),
    .Z(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11235_ (.I(_05442_),
    .Z(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11236_ (.A1(_04223_),
    .A2(_05527_),
    .ZN(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11237_ (.I(_05528_),
    .Z(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11238_ (.I0(_05500_),
    .I1(\u2.mem[152][0] ),
    .S(_05529_),
    .Z(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11239_ (.I(_05530_),
    .Z(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11240_ (.I0(_05505_),
    .I1(\u2.mem[152][1] ),
    .S(_05529_),
    .Z(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11241_ (.I(_05531_),
    .Z(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11242_ (.I0(_05508_),
    .I1(\u2.mem[152][2] ),
    .S(_05529_),
    .Z(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11243_ (.I(_05532_),
    .Z(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11244_ (.I0(_05511_),
    .I1(\u2.mem[152][3] ),
    .S(_05529_),
    .Z(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11245_ (.I(_05533_),
    .Z(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11246_ (.I0(_05514_),
    .I1(\u2.mem[152][4] ),
    .S(_05528_),
    .Z(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11247_ (.I(_05534_),
    .Z(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11248_ (.I0(_05517_),
    .I1(\u2.mem[152][5] ),
    .S(_05528_),
    .Z(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11249_ (.I(_05535_),
    .Z(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11250_ (.A1(_04248_),
    .A2(_05527_),
    .ZN(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11251_ (.I(_05536_),
    .Z(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11252_ (.I0(_05500_),
    .I1(\u2.mem[153][0] ),
    .S(_05537_),
    .Z(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11253_ (.I(_05538_),
    .Z(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11254_ (.I0(_05505_),
    .I1(\u2.mem[153][1] ),
    .S(_05537_),
    .Z(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11255_ (.I(_05539_),
    .Z(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11256_ (.I0(_05508_),
    .I1(\u2.mem[153][2] ),
    .S(_05537_),
    .Z(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11257_ (.I(_05540_),
    .Z(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11258_ (.I0(_05511_),
    .I1(\u2.mem[153][3] ),
    .S(_05537_),
    .Z(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11259_ (.I(_05541_),
    .Z(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11260_ (.I0(_05514_),
    .I1(\u2.mem[153][4] ),
    .S(_05536_),
    .Z(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11261_ (.I(_05542_),
    .Z(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11262_ (.I0(_05517_),
    .I1(\u2.mem[153][5] ),
    .S(_05536_),
    .Z(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11263_ (.I(_05543_),
    .Z(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11264_ (.I(_05499_),
    .Z(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11265_ (.A1(_04287_),
    .A2(_05527_),
    .ZN(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11266_ (.I(_05545_),
    .Z(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11267_ (.I0(_05544_),
    .I1(\u2.mem[154][0] ),
    .S(_05546_),
    .Z(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11268_ (.I(_05547_),
    .Z(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11269_ (.I(_05504_),
    .Z(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11270_ (.I0(_05548_),
    .I1(\u2.mem[154][1] ),
    .S(_05546_),
    .Z(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11271_ (.I(_05549_),
    .Z(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11272_ (.I(_05507_),
    .Z(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11273_ (.I0(_05550_),
    .I1(\u2.mem[154][2] ),
    .S(_05546_),
    .Z(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11274_ (.I(_05551_),
    .Z(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11275_ (.I(_05510_),
    .Z(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11276_ (.I0(_05552_),
    .I1(\u2.mem[154][3] ),
    .S(_05546_),
    .Z(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11277_ (.I(_05553_),
    .Z(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11278_ (.I(_05513_),
    .Z(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11279_ (.I0(_05554_),
    .I1(\u2.mem[154][4] ),
    .S(_05545_),
    .Z(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11280_ (.I(_05555_),
    .Z(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11281_ (.I(_05516_),
    .Z(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11282_ (.I0(_05556_),
    .I1(\u2.mem[154][5] ),
    .S(_05545_),
    .Z(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11283_ (.I(_05557_),
    .Z(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11284_ (.A1(_04310_),
    .A2(_05527_),
    .ZN(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11285_ (.I(_05558_),
    .Z(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11286_ (.I0(_05544_),
    .I1(\u2.mem[155][0] ),
    .S(_05559_),
    .Z(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11287_ (.I(_05560_),
    .Z(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11288_ (.I0(_05548_),
    .I1(\u2.mem[155][1] ),
    .S(_05559_),
    .Z(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11289_ (.I(_05561_),
    .Z(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11290_ (.I0(_05550_),
    .I1(\u2.mem[155][2] ),
    .S(_05559_),
    .Z(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11291_ (.I(_05562_),
    .Z(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11292_ (.I0(_05552_),
    .I1(\u2.mem[155][3] ),
    .S(_05559_),
    .Z(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11293_ (.I(_05563_),
    .Z(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11294_ (.I0(_05554_),
    .I1(\u2.mem[155][4] ),
    .S(_05558_),
    .Z(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11295_ (.I(_05564_),
    .Z(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11296_ (.I0(_05556_),
    .I1(\u2.mem[155][5] ),
    .S(_05558_),
    .Z(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11297_ (.I(_05565_),
    .Z(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11298_ (.I(_05442_),
    .Z(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11299_ (.A1(_04333_),
    .A2(_05566_),
    .ZN(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11300_ (.I(_05567_),
    .Z(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11301_ (.I0(_05544_),
    .I1(\u2.mem[156][0] ),
    .S(_05568_),
    .Z(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11302_ (.I(_05569_),
    .Z(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11303_ (.I0(_05548_),
    .I1(\u2.mem[156][1] ),
    .S(_05568_),
    .Z(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11304_ (.I(_05570_),
    .Z(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11305_ (.I0(_05550_),
    .I1(\u2.mem[156][2] ),
    .S(_05568_),
    .Z(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11306_ (.I(_05571_),
    .Z(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11307_ (.I0(_05552_),
    .I1(\u2.mem[156][3] ),
    .S(_05568_),
    .Z(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11308_ (.I(_05572_),
    .Z(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11309_ (.I0(_05554_),
    .I1(\u2.mem[156][4] ),
    .S(_05567_),
    .Z(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11310_ (.I(_05573_),
    .Z(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11311_ (.I0(_05556_),
    .I1(\u2.mem[156][5] ),
    .S(_05567_),
    .Z(_05574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11312_ (.I(_05574_),
    .Z(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11313_ (.A1(_05411_),
    .A2(_05566_),
    .ZN(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11314_ (.I(_05575_),
    .Z(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11315_ (.I0(_05544_),
    .I1(\u2.mem[157][0] ),
    .S(_05576_),
    .Z(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11316_ (.I(_05577_),
    .Z(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11317_ (.I0(_05548_),
    .I1(\u2.mem[157][1] ),
    .S(_05576_),
    .Z(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11318_ (.I(_05578_),
    .Z(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11319_ (.I0(_05550_),
    .I1(\u2.mem[157][2] ),
    .S(_05576_),
    .Z(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11320_ (.I(_05579_),
    .Z(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11321_ (.I0(_05552_),
    .I1(\u2.mem[157][3] ),
    .S(_05576_),
    .Z(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11322_ (.I(_05580_),
    .Z(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11323_ (.I0(_05554_),
    .I1(\u2.mem[157][4] ),
    .S(_05575_),
    .Z(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11324_ (.I(_05581_),
    .Z(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11325_ (.I0(_05556_),
    .I1(\u2.mem[157][5] ),
    .S(_05575_),
    .Z(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11326_ (.I(_05582_),
    .Z(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11327_ (.I(_05499_),
    .Z(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11328_ (.A1(_04393_),
    .A2(_05566_),
    .ZN(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11329_ (.I(_05584_),
    .Z(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11330_ (.I0(_05583_),
    .I1(\u2.mem[158][0] ),
    .S(_05585_),
    .Z(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11331_ (.I(_05586_),
    .Z(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11332_ (.I(_05504_),
    .Z(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11333_ (.I0(_05587_),
    .I1(\u2.mem[158][1] ),
    .S(_05585_),
    .Z(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11334_ (.I(_05588_),
    .Z(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11335_ (.I(_05507_),
    .Z(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11336_ (.I0(_05589_),
    .I1(\u2.mem[158][2] ),
    .S(_05585_),
    .Z(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11337_ (.I(_05590_),
    .Z(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11338_ (.I(_05510_),
    .Z(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11339_ (.I0(_05591_),
    .I1(\u2.mem[158][3] ),
    .S(_05585_),
    .Z(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11340_ (.I(_05592_),
    .Z(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11341_ (.I(_05513_),
    .Z(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11342_ (.I0(_05593_),
    .I1(\u2.mem[158][4] ),
    .S(_05584_),
    .Z(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11343_ (.I(_05594_),
    .Z(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11344_ (.I(_05516_),
    .Z(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11345_ (.I0(_05595_),
    .I1(\u2.mem[158][5] ),
    .S(_05584_),
    .Z(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11346_ (.I(_05596_),
    .Z(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11347_ (.A1(_04417_),
    .A2(_05566_),
    .ZN(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11348_ (.I(_05597_),
    .Z(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11349_ (.I0(_05583_),
    .I1(\u2.mem[159][0] ),
    .S(_05598_),
    .Z(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11350_ (.I(_05599_),
    .Z(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11351_ (.I0(_05587_),
    .I1(\u2.mem[159][1] ),
    .S(_05598_),
    .Z(_05600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11352_ (.I(_05600_),
    .Z(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11353_ (.I0(_05589_),
    .I1(\u2.mem[159][2] ),
    .S(_05598_),
    .Z(_05601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11354_ (.I(_05601_),
    .Z(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11355_ (.I0(_05591_),
    .I1(\u2.mem[159][3] ),
    .S(_05598_),
    .Z(_05602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11356_ (.I(_05602_),
    .Z(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11357_ (.I0(_05593_),
    .I1(\u2.mem[159][4] ),
    .S(_05597_),
    .Z(_05603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11358_ (.I(_05603_),
    .Z(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11359_ (.I0(_05595_),
    .I1(\u2.mem[159][5] ),
    .S(_05597_),
    .Z(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11360_ (.I(_05604_),
    .Z(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11361_ (.A1(_04439_),
    .A2(_05274_),
    .ZN(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11362_ (.I(_05605_),
    .Z(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11363_ (.A1(_03487_),
    .A2(_05606_),
    .ZN(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11364_ (.I(_05607_),
    .Z(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11365_ (.I0(_05583_),
    .I1(\u2.mem[160][0] ),
    .S(_05608_),
    .Z(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11366_ (.I(_05609_),
    .Z(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11367_ (.I0(_05587_),
    .I1(\u2.mem[160][1] ),
    .S(_05608_),
    .Z(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11368_ (.I(_05610_),
    .Z(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11369_ (.I0(_05589_),
    .I1(\u2.mem[160][2] ),
    .S(_05608_),
    .Z(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11370_ (.I(_05611_),
    .Z(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11371_ (.I0(_05591_),
    .I1(\u2.mem[160][3] ),
    .S(_05608_),
    .Z(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11372_ (.I(_05612_),
    .Z(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11373_ (.I0(_05593_),
    .I1(\u2.mem[160][4] ),
    .S(_05607_),
    .Z(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11374_ (.I(_05613_),
    .Z(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11375_ (.I0(_05595_),
    .I1(\u2.mem[160][5] ),
    .S(_05607_),
    .Z(_05614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11376_ (.I(_05614_),
    .Z(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11377_ (.A1(_05285_),
    .A2(_05606_),
    .ZN(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11378_ (.I(_05615_),
    .Z(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11379_ (.I0(_05583_),
    .I1(\u2.mem[161][0] ),
    .S(_05616_),
    .Z(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11380_ (.I(_05617_),
    .Z(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11381_ (.I0(_05587_),
    .I1(\u2.mem[161][1] ),
    .S(_05616_),
    .Z(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11382_ (.I(_05618_),
    .Z(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11383_ (.I0(_05589_),
    .I1(\u2.mem[161][2] ),
    .S(_05616_),
    .Z(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11384_ (.I(_05619_),
    .Z(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11385_ (.I0(_05591_),
    .I1(\u2.mem[161][3] ),
    .S(_05616_),
    .Z(_05620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11386_ (.I(_05620_),
    .Z(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11387_ (.I0(_05593_),
    .I1(\u2.mem[161][4] ),
    .S(_05615_),
    .Z(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11388_ (.I(_05621_),
    .Z(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11389_ (.I0(_05595_),
    .I1(\u2.mem[161][5] ),
    .S(_05615_),
    .Z(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11390_ (.I(_05622_),
    .Z(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11391_ (.I(_05499_),
    .Z(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11392_ (.A1(_05295_),
    .A2(_05606_),
    .ZN(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11393_ (.I(_05624_),
    .Z(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11394_ (.I0(_05623_),
    .I1(\u2.mem[162][0] ),
    .S(_05625_),
    .Z(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11395_ (.I(_05626_),
    .Z(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11396_ (.I(_05504_),
    .Z(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11397_ (.I0(_05627_),
    .I1(\u2.mem[162][1] ),
    .S(_05625_),
    .Z(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11398_ (.I(_05628_),
    .Z(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11399_ (.I(_05507_),
    .Z(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11400_ (.I0(_05629_),
    .I1(\u2.mem[162][2] ),
    .S(_05625_),
    .Z(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11401_ (.I(_05630_),
    .Z(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11402_ (.I(_05510_),
    .Z(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11403_ (.I0(_05631_),
    .I1(\u2.mem[162][3] ),
    .S(_05625_),
    .Z(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11404_ (.I(_05632_),
    .Z(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11405_ (.I(_05513_),
    .Z(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11406_ (.I0(_05633_),
    .I1(\u2.mem[162][4] ),
    .S(_05624_),
    .Z(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11407_ (.I(_05634_),
    .Z(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11408_ (.I(_05516_),
    .Z(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11409_ (.I0(_05635_),
    .I1(\u2.mem[162][5] ),
    .S(_05624_),
    .Z(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11410_ (.I(_05636_),
    .Z(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11411_ (.A1(_04071_),
    .A2(_05606_),
    .ZN(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11412_ (.I(_05637_),
    .Z(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11413_ (.I0(_05623_),
    .I1(\u2.mem[163][0] ),
    .S(_05638_),
    .Z(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11414_ (.I(_05639_),
    .Z(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11415_ (.I0(_05627_),
    .I1(\u2.mem[163][1] ),
    .S(_05638_),
    .Z(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11416_ (.I(_05640_),
    .Z(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11417_ (.I0(_05629_),
    .I1(\u2.mem[163][2] ),
    .S(_05638_),
    .Z(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11418_ (.I(_05641_),
    .Z(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11419_ (.I0(_05631_),
    .I1(\u2.mem[163][3] ),
    .S(_05638_),
    .Z(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11420_ (.I(_05642_),
    .Z(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11421_ (.I0(_05633_),
    .I1(\u2.mem[163][4] ),
    .S(_05637_),
    .Z(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11422_ (.I(_05643_),
    .Z(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11423_ (.I0(_05635_),
    .I1(\u2.mem[163][5] ),
    .S(_05637_),
    .Z(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11424_ (.I(_05644_),
    .Z(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11425_ (.I(_05605_),
    .Z(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11426_ (.A1(_04094_),
    .A2(_05645_),
    .ZN(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11427_ (.I(_05646_),
    .Z(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11428_ (.I0(_05623_),
    .I1(\u2.mem[164][0] ),
    .S(_05647_),
    .Z(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11429_ (.I(_05648_),
    .Z(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11430_ (.I0(_05627_),
    .I1(\u2.mem[164][1] ),
    .S(_05647_),
    .Z(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11431_ (.I(_05649_),
    .Z(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11432_ (.I0(_05629_),
    .I1(\u2.mem[164][2] ),
    .S(_05647_),
    .Z(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11433_ (.I(_05650_),
    .Z(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11434_ (.I0(_05631_),
    .I1(\u2.mem[164][3] ),
    .S(_05647_),
    .Z(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11435_ (.I(_05651_),
    .Z(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11436_ (.I0(_05633_),
    .I1(\u2.mem[164][4] ),
    .S(_05646_),
    .Z(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11437_ (.I(_05652_),
    .Z(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11438_ (.I0(_05635_),
    .I1(\u2.mem[164][5] ),
    .S(_05646_),
    .Z(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11439_ (.I(_05653_),
    .Z(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11440_ (.A1(_04120_),
    .A2(_05645_),
    .ZN(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11441_ (.I(_05654_),
    .Z(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11442_ (.I0(_05623_),
    .I1(\u2.mem[165][0] ),
    .S(_05655_),
    .Z(_05656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11443_ (.I(_05656_),
    .Z(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11444_ (.I0(_05627_),
    .I1(\u2.mem[165][1] ),
    .S(_05655_),
    .Z(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11445_ (.I(_05657_),
    .Z(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11446_ (.I0(_05629_),
    .I1(\u2.mem[165][2] ),
    .S(_05655_),
    .Z(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11447_ (.I(_05658_),
    .Z(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11448_ (.I0(_05631_),
    .I1(\u2.mem[165][3] ),
    .S(_05655_),
    .Z(_05659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11449_ (.I(_05659_),
    .Z(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11450_ (.I0(_05633_),
    .I1(\u2.mem[165][4] ),
    .S(_05654_),
    .Z(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11451_ (.I(_05660_),
    .Z(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11452_ (.I0(_05635_),
    .I1(\u2.mem[165][5] ),
    .S(_05654_),
    .Z(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11453_ (.I(_05661_),
    .Z(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11454_ (.I(_03491_),
    .Z(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11455_ (.I(_05662_),
    .Z(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11456_ (.A1(_04179_),
    .A2(_05645_),
    .ZN(_05664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11457_ (.I(_05664_),
    .Z(_05665_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11458_ (.I0(_05663_),
    .I1(\u2.mem[166][0] ),
    .S(_05665_),
    .Z(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11459_ (.I(_05666_),
    .Z(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11460_ (.I(_03496_),
    .Z(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11461_ (.I(_05667_),
    .Z(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11462_ (.I0(_05668_),
    .I1(\u2.mem[166][1] ),
    .S(_05665_),
    .Z(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11463_ (.I(_05669_),
    .Z(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11464_ (.I(_03499_),
    .Z(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11465_ (.I(_05670_),
    .Z(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11466_ (.I0(_05671_),
    .I1(\u2.mem[166][2] ),
    .S(_05665_),
    .Z(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11467_ (.I(_05672_),
    .Z(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11468_ (.I(_03502_),
    .Z(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11469_ (.I(_05673_),
    .Z(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11470_ (.I0(_05674_),
    .I1(\u2.mem[166][3] ),
    .S(_05665_),
    .Z(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11471_ (.I(_05675_),
    .Z(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11472_ (.I(_03506_),
    .Z(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11473_ (.I(_05676_),
    .Z(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11474_ (.I0(_05677_),
    .I1(\u2.mem[166][4] ),
    .S(_05664_),
    .Z(_05678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11475_ (.I(_05678_),
    .Z(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11476_ (.I(_03510_),
    .Z(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11477_ (.I(_05679_),
    .Z(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11478_ (.I0(_05680_),
    .I1(\u2.mem[166][5] ),
    .S(_05664_),
    .Z(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11479_ (.I(_05681_),
    .Z(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11480_ (.A1(_05354_),
    .A2(_05645_),
    .ZN(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11481_ (.I(_05682_),
    .Z(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11482_ (.I0(_05663_),
    .I1(\u2.mem[167][0] ),
    .S(_05683_),
    .Z(_05684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11483_ (.I(_05684_),
    .Z(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11484_ (.I0(_05668_),
    .I1(\u2.mem[167][1] ),
    .S(_05683_),
    .Z(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11485_ (.I(_05685_),
    .Z(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11486_ (.I0(_05671_),
    .I1(\u2.mem[167][2] ),
    .S(_05683_),
    .Z(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11487_ (.I(_05686_),
    .Z(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11488_ (.I0(_05674_),
    .I1(\u2.mem[167][3] ),
    .S(_05683_),
    .Z(_05687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11489_ (.I(_05687_),
    .Z(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11490_ (.I0(_05677_),
    .I1(\u2.mem[167][4] ),
    .S(_05682_),
    .Z(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11491_ (.I(_05688_),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11492_ (.I0(_05680_),
    .I1(\u2.mem[167][5] ),
    .S(_05682_),
    .Z(_05689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11493_ (.I(_05689_),
    .Z(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11494_ (.I(_05605_),
    .Z(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11495_ (.A1(_04223_),
    .A2(_05690_),
    .ZN(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11496_ (.I(_05691_),
    .Z(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11497_ (.I0(_05663_),
    .I1(\u2.mem[168][0] ),
    .S(_05692_),
    .Z(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11498_ (.I(_05693_),
    .Z(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11499_ (.I0(_05668_),
    .I1(\u2.mem[168][1] ),
    .S(_05692_),
    .Z(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11500_ (.I(_05694_),
    .Z(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11501_ (.I0(_05671_),
    .I1(\u2.mem[168][2] ),
    .S(_05692_),
    .Z(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11502_ (.I(_05695_),
    .Z(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11503_ (.I0(_05674_),
    .I1(\u2.mem[168][3] ),
    .S(_05692_),
    .Z(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11504_ (.I(_05696_),
    .Z(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11505_ (.I0(_05677_),
    .I1(\u2.mem[168][4] ),
    .S(_05691_),
    .Z(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11506_ (.I(_05697_),
    .Z(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11507_ (.I0(_05680_),
    .I1(\u2.mem[168][5] ),
    .S(_05691_),
    .Z(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11508_ (.I(_05698_),
    .Z(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11509_ (.A1(_04248_),
    .A2(_05690_),
    .ZN(_05699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11510_ (.I(_05699_),
    .Z(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11511_ (.I0(_05663_),
    .I1(\u2.mem[169][0] ),
    .S(_05700_),
    .Z(_05701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11512_ (.I(_05701_),
    .Z(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11513_ (.I0(_05668_),
    .I1(\u2.mem[169][1] ),
    .S(_05700_),
    .Z(_05702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11514_ (.I(_05702_),
    .Z(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11515_ (.I0(_05671_),
    .I1(\u2.mem[169][2] ),
    .S(_05700_),
    .Z(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11516_ (.I(_05703_),
    .Z(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11517_ (.I0(_05674_),
    .I1(\u2.mem[169][3] ),
    .S(_05700_),
    .Z(_05704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11518_ (.I(_05704_),
    .Z(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11519_ (.I0(_05677_),
    .I1(\u2.mem[169][4] ),
    .S(_05699_),
    .Z(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11520_ (.I(_05705_),
    .Z(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11521_ (.I0(_05680_),
    .I1(\u2.mem[169][5] ),
    .S(_05699_),
    .Z(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11522_ (.I(_05706_),
    .Z(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11523_ (.I(_05662_),
    .Z(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11524_ (.A1(_04287_),
    .A2(_05690_),
    .ZN(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11525_ (.I(_05708_),
    .Z(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11526_ (.I0(_05707_),
    .I1(\u2.mem[170][0] ),
    .S(_05709_),
    .Z(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11527_ (.I(_05710_),
    .Z(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11528_ (.I(_05667_),
    .Z(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11529_ (.I0(_05711_),
    .I1(\u2.mem[170][1] ),
    .S(_05709_),
    .Z(_05712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11530_ (.I(_05712_),
    .Z(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11531_ (.I(_05670_),
    .Z(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11532_ (.I0(_05713_),
    .I1(\u2.mem[170][2] ),
    .S(_05709_),
    .Z(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11533_ (.I(_05714_),
    .Z(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11534_ (.I(_05673_),
    .Z(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11535_ (.I0(_05715_),
    .I1(\u2.mem[170][3] ),
    .S(_05709_),
    .Z(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11536_ (.I(_05716_),
    .Z(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11537_ (.I(_05676_),
    .Z(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11538_ (.I0(_05717_),
    .I1(\u2.mem[170][4] ),
    .S(_05708_),
    .Z(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11539_ (.I(_05718_),
    .Z(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11540_ (.I(_05679_),
    .Z(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11541_ (.I0(_05719_),
    .I1(\u2.mem[170][5] ),
    .S(_05708_),
    .Z(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11542_ (.I(_05720_),
    .Z(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11543_ (.A1(_04310_),
    .A2(_05690_),
    .ZN(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11544_ (.I(_05721_),
    .Z(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11545_ (.I0(_05707_),
    .I1(\u2.mem[171][0] ),
    .S(_05722_),
    .Z(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11546_ (.I(_05723_),
    .Z(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11547_ (.I0(_05711_),
    .I1(\u2.mem[171][1] ),
    .S(_05722_),
    .Z(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11548_ (.I(_05724_),
    .Z(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11549_ (.I0(_05713_),
    .I1(\u2.mem[171][2] ),
    .S(_05722_),
    .Z(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11550_ (.I(_05725_),
    .Z(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11551_ (.I0(_05715_),
    .I1(\u2.mem[171][3] ),
    .S(_05722_),
    .Z(_05726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11552_ (.I(_05726_),
    .Z(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11553_ (.I0(_05717_),
    .I1(\u2.mem[171][4] ),
    .S(_05721_),
    .Z(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11554_ (.I(_05727_),
    .Z(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11555_ (.I0(_05719_),
    .I1(\u2.mem[171][5] ),
    .S(_05721_),
    .Z(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11556_ (.I(_05728_),
    .Z(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11557_ (.I(_05605_),
    .Z(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11558_ (.A1(_04333_),
    .A2(_05729_),
    .ZN(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11559_ (.I(_05730_),
    .Z(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11560_ (.I0(_05707_),
    .I1(\u2.mem[172][0] ),
    .S(_05731_),
    .Z(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11561_ (.I(_05732_),
    .Z(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11562_ (.I0(_05711_),
    .I1(\u2.mem[172][1] ),
    .S(_05731_),
    .Z(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11563_ (.I(_05733_),
    .Z(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11564_ (.I0(_05713_),
    .I1(\u2.mem[172][2] ),
    .S(_05731_),
    .Z(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11565_ (.I(_05734_),
    .Z(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11566_ (.I0(_05715_),
    .I1(\u2.mem[172][3] ),
    .S(_05731_),
    .Z(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11567_ (.I(_05735_),
    .Z(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11568_ (.I0(_05717_),
    .I1(\u2.mem[172][4] ),
    .S(_05730_),
    .Z(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11569_ (.I(_05736_),
    .Z(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11570_ (.I0(_05719_),
    .I1(\u2.mem[172][5] ),
    .S(_05730_),
    .Z(_05737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11571_ (.I(_05737_),
    .Z(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11572_ (.A1(_05411_),
    .A2(_05729_),
    .ZN(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11573_ (.I(_05738_),
    .Z(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11574_ (.I0(_05707_),
    .I1(\u2.mem[173][0] ),
    .S(_05739_),
    .Z(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11575_ (.I(_05740_),
    .Z(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11576_ (.I0(_05711_),
    .I1(\u2.mem[173][1] ),
    .S(_05739_),
    .Z(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11577_ (.I(_05741_),
    .Z(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11578_ (.I0(_05713_),
    .I1(\u2.mem[173][2] ),
    .S(_05739_),
    .Z(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11579_ (.I(_05742_),
    .Z(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11580_ (.I0(_05715_),
    .I1(\u2.mem[173][3] ),
    .S(_05739_),
    .Z(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11581_ (.I(_05743_),
    .Z(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11582_ (.I0(_05717_),
    .I1(\u2.mem[173][4] ),
    .S(_05738_),
    .Z(_05744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11583_ (.I(_05744_),
    .Z(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11584_ (.I0(_05719_),
    .I1(\u2.mem[173][5] ),
    .S(_05738_),
    .Z(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11585_ (.I(_05745_),
    .Z(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11586_ (.I(_05662_),
    .Z(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11587_ (.A1(_04393_),
    .A2(_05729_),
    .ZN(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11588_ (.I(_05747_),
    .Z(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11589_ (.I0(_05746_),
    .I1(\u2.mem[174][0] ),
    .S(_05748_),
    .Z(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11590_ (.I(_05749_),
    .Z(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11591_ (.I(_05667_),
    .Z(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11592_ (.I0(_05750_),
    .I1(\u2.mem[174][1] ),
    .S(_05748_),
    .Z(_05751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11593_ (.I(_05751_),
    .Z(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11594_ (.I(_05670_),
    .Z(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11595_ (.I0(_05752_),
    .I1(\u2.mem[174][2] ),
    .S(_05748_),
    .Z(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11596_ (.I(_05753_),
    .Z(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11597_ (.I(_05673_),
    .Z(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11598_ (.I0(_05754_),
    .I1(\u2.mem[174][3] ),
    .S(_05748_),
    .Z(_05755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11599_ (.I(_05755_),
    .Z(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11600_ (.I(_05676_),
    .Z(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11601_ (.I0(_05756_),
    .I1(\u2.mem[174][4] ),
    .S(_05747_),
    .Z(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11602_ (.I(_05757_),
    .Z(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11603_ (.I(_05679_),
    .Z(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11604_ (.I0(_05758_),
    .I1(\u2.mem[174][5] ),
    .S(_05747_),
    .Z(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11605_ (.I(_05759_),
    .Z(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11606_ (.A1(_04416_),
    .A2(_05729_),
    .ZN(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11607_ (.I(_05760_),
    .Z(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11608_ (.I0(_05746_),
    .I1(\u2.mem[175][0] ),
    .S(_05761_),
    .Z(_05762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11609_ (.I(_05762_),
    .Z(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11610_ (.I0(_05750_),
    .I1(\u2.mem[175][1] ),
    .S(_05761_),
    .Z(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11611_ (.I(_05763_),
    .Z(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11612_ (.I0(_05752_),
    .I1(\u2.mem[175][2] ),
    .S(_05761_),
    .Z(_05764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11613_ (.I(_05764_),
    .Z(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11614_ (.I0(_05754_),
    .I1(\u2.mem[175][3] ),
    .S(_05761_),
    .Z(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11615_ (.I(_05765_),
    .Z(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11616_ (.I0(_05756_),
    .I1(\u2.mem[175][4] ),
    .S(_05760_),
    .Z(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11617_ (.I(_05766_),
    .Z(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11618_ (.I0(_05758_),
    .I1(\u2.mem[175][5] ),
    .S(_05760_),
    .Z(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11619_ (.I(_05767_),
    .Z(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11620_ (.A1(_04861_),
    .A2(_05274_),
    .ZN(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11621_ (.I(_05768_),
    .Z(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11622_ (.A1(_03487_),
    .A2(_05769_),
    .ZN(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11623_ (.I(_05770_),
    .Z(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11624_ (.I0(_05746_),
    .I1(\u2.mem[176][0] ),
    .S(_05771_),
    .Z(_05772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11625_ (.I(_05772_),
    .Z(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11626_ (.I0(_05750_),
    .I1(\u2.mem[176][1] ),
    .S(_05771_),
    .Z(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11627_ (.I(_05773_),
    .Z(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11628_ (.I0(_05752_),
    .I1(\u2.mem[176][2] ),
    .S(_05771_),
    .Z(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11629_ (.I(_05774_),
    .Z(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11630_ (.I0(_05754_),
    .I1(\u2.mem[176][3] ),
    .S(_05771_),
    .Z(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11631_ (.I(_05775_),
    .Z(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11632_ (.I0(_05756_),
    .I1(\u2.mem[176][4] ),
    .S(_05770_),
    .Z(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11633_ (.I(_05776_),
    .Z(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11634_ (.I0(_05758_),
    .I1(\u2.mem[176][5] ),
    .S(_05770_),
    .Z(_05777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11635_ (.I(_05777_),
    .Z(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11636_ (.A1(_05285_),
    .A2(_05769_),
    .ZN(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11637_ (.I(_05778_),
    .Z(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11638_ (.I0(_05746_),
    .I1(\u2.mem[177][0] ),
    .S(_05779_),
    .Z(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11639_ (.I(_05780_),
    .Z(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11640_ (.I0(_05750_),
    .I1(\u2.mem[177][1] ),
    .S(_05779_),
    .Z(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11641_ (.I(_05781_),
    .Z(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11642_ (.I0(_05752_),
    .I1(\u2.mem[177][2] ),
    .S(_05779_),
    .Z(_05782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11643_ (.I(_05782_),
    .Z(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11644_ (.I0(_05754_),
    .I1(\u2.mem[177][3] ),
    .S(_05779_),
    .Z(_05783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11645_ (.I(_05783_),
    .Z(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11646_ (.I0(_05756_),
    .I1(\u2.mem[177][4] ),
    .S(_05778_),
    .Z(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11647_ (.I(_05784_),
    .Z(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11648_ (.I0(_05758_),
    .I1(\u2.mem[177][5] ),
    .S(_05778_),
    .Z(_05785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11649_ (.I(_05785_),
    .Z(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11650_ (.I(_05662_),
    .Z(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11651_ (.A1(_05295_),
    .A2(_05769_),
    .ZN(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11652_ (.I(_05787_),
    .Z(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11653_ (.I0(_05786_),
    .I1(\u2.mem[178][0] ),
    .S(_05788_),
    .Z(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11654_ (.I(_05789_),
    .Z(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11655_ (.I(_05667_),
    .Z(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11656_ (.I0(_05790_),
    .I1(\u2.mem[178][1] ),
    .S(_05788_),
    .Z(_05791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11657_ (.I(_05791_),
    .Z(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11658_ (.I(_05670_),
    .Z(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11659_ (.I0(_05792_),
    .I1(\u2.mem[178][2] ),
    .S(_05788_),
    .Z(_05793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11660_ (.I(_05793_),
    .Z(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11661_ (.I(_05673_),
    .Z(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11662_ (.I0(_05794_),
    .I1(\u2.mem[178][3] ),
    .S(_05788_),
    .Z(_05795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11663_ (.I(_05795_),
    .Z(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11664_ (.I(_05676_),
    .Z(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11665_ (.I0(_05796_),
    .I1(\u2.mem[178][4] ),
    .S(_05787_),
    .Z(_05797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11666_ (.I(_05797_),
    .Z(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11667_ (.I(_05679_),
    .Z(_05798_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11668_ (.I0(_05798_),
    .I1(\u2.mem[178][5] ),
    .S(_05787_),
    .Z(_05799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11669_ (.I(_05799_),
    .Z(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11670_ (.A1(_04071_),
    .A2(_05769_),
    .ZN(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11671_ (.I(_05800_),
    .Z(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11672_ (.I0(_05786_),
    .I1(\u2.mem[179][0] ),
    .S(_05801_),
    .Z(_05802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11673_ (.I(_05802_),
    .Z(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11674_ (.I0(_05790_),
    .I1(\u2.mem[179][1] ),
    .S(_05801_),
    .Z(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11675_ (.I(_05803_),
    .Z(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11676_ (.I0(_05792_),
    .I1(\u2.mem[179][2] ),
    .S(_05801_),
    .Z(_05804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11677_ (.I(_05804_),
    .Z(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11678_ (.I0(_05794_),
    .I1(\u2.mem[179][3] ),
    .S(_05801_),
    .Z(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11679_ (.I(_05805_),
    .Z(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11680_ (.I0(_05796_),
    .I1(\u2.mem[179][4] ),
    .S(_05800_),
    .Z(_05806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11681_ (.I(_05806_),
    .Z(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11682_ (.I0(_05798_),
    .I1(\u2.mem[179][5] ),
    .S(_05800_),
    .Z(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11683_ (.I(_05807_),
    .Z(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11684_ (.I(_05768_),
    .Z(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11685_ (.A1(_04094_),
    .A2(_05808_),
    .ZN(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11686_ (.I(_05809_),
    .Z(_05810_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11687_ (.I0(_05786_),
    .I1(\u2.mem[180][0] ),
    .S(_05810_),
    .Z(_05811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11688_ (.I(_05811_),
    .Z(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11689_ (.I0(_05790_),
    .I1(\u2.mem[180][1] ),
    .S(_05810_),
    .Z(_05812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11690_ (.I(_05812_),
    .Z(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11691_ (.I0(_05792_),
    .I1(\u2.mem[180][2] ),
    .S(_05810_),
    .Z(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11692_ (.I(_05813_),
    .Z(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11693_ (.I0(_05794_),
    .I1(\u2.mem[180][3] ),
    .S(_05810_),
    .Z(_05814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11694_ (.I(_05814_),
    .Z(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11695_ (.I0(_05796_),
    .I1(\u2.mem[180][4] ),
    .S(_05809_),
    .Z(_05815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11696_ (.I(_05815_),
    .Z(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11697_ (.I0(_05798_),
    .I1(\u2.mem[180][5] ),
    .S(_05809_),
    .Z(_05816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11698_ (.I(_05816_),
    .Z(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11699_ (.A1(_04120_),
    .A2(_05808_),
    .ZN(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11700_ (.I(_05817_),
    .Z(_05818_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11701_ (.I0(_05786_),
    .I1(\u2.mem[181][0] ),
    .S(_05818_),
    .Z(_05819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11702_ (.I(_05819_),
    .Z(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11703_ (.I0(_05790_),
    .I1(\u2.mem[181][1] ),
    .S(_05818_),
    .Z(_05820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11704_ (.I(_05820_),
    .Z(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11705_ (.I0(_05792_),
    .I1(\u2.mem[181][2] ),
    .S(_05818_),
    .Z(_05821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11706_ (.I(_05821_),
    .Z(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11707_ (.I0(_05794_),
    .I1(\u2.mem[181][3] ),
    .S(_05818_),
    .Z(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11708_ (.I(_05822_),
    .Z(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11709_ (.I0(_05796_),
    .I1(\u2.mem[181][4] ),
    .S(_05817_),
    .Z(_05823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11710_ (.I(_05823_),
    .Z(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11711_ (.I0(_05798_),
    .I1(\u2.mem[181][5] ),
    .S(_05817_),
    .Z(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11712_ (.I(_05824_),
    .Z(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11713_ (.I(_03655_),
    .Z(_05825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11714_ (.A1(_04179_),
    .A2(_05808_),
    .ZN(_05826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11715_ (.I(_05826_),
    .Z(_05827_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11716_ (.I0(_05825_),
    .I1(\u2.mem[182][0] ),
    .S(_05827_),
    .Z(_05828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11717_ (.I(_05828_),
    .Z(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11718_ (.I(_03662_),
    .Z(_05829_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11719_ (.I0(_05829_),
    .I1(\u2.mem[182][1] ),
    .S(_05827_),
    .Z(_05830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11720_ (.I(_05830_),
    .Z(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11721_ (.I(_03666_),
    .Z(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11722_ (.I0(_05831_),
    .I1(\u2.mem[182][2] ),
    .S(_05827_),
    .Z(_05832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11723_ (.I(_05832_),
    .Z(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11724_ (.I(_03670_),
    .Z(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11725_ (.I0(_05833_),
    .I1(\u2.mem[182][3] ),
    .S(_05827_),
    .Z(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11726_ (.I(_05834_),
    .Z(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11727_ (.I(_03674_),
    .Z(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11728_ (.I0(_05835_),
    .I1(\u2.mem[182][4] ),
    .S(_05826_),
    .Z(_05836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11729_ (.I(_05836_),
    .Z(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11730_ (.I(_03679_),
    .Z(_05837_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11731_ (.I0(_05837_),
    .I1(\u2.mem[182][5] ),
    .S(_05826_),
    .Z(_05838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11732_ (.I(_05838_),
    .Z(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11733_ (.A1(_05354_),
    .A2(_05808_),
    .ZN(_05839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11734_ (.I(_05839_),
    .Z(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11735_ (.I0(_05825_),
    .I1(\u2.mem[183][0] ),
    .S(_05840_),
    .Z(_05841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11736_ (.I(_05841_),
    .Z(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11737_ (.I0(_05829_),
    .I1(\u2.mem[183][1] ),
    .S(_05840_),
    .Z(_05842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11738_ (.I(_05842_),
    .Z(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11739_ (.I0(_05831_),
    .I1(\u2.mem[183][2] ),
    .S(_05840_),
    .Z(_05843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11740_ (.I(_05843_),
    .Z(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11741_ (.I0(_05833_),
    .I1(\u2.mem[183][3] ),
    .S(_05840_),
    .Z(_05844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11742_ (.I(_05844_),
    .Z(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11743_ (.I0(_05835_),
    .I1(\u2.mem[183][4] ),
    .S(_05839_),
    .Z(_05845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11744_ (.I(_05845_),
    .Z(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11745_ (.I0(_05837_),
    .I1(\u2.mem[183][5] ),
    .S(_05839_),
    .Z(_05846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11746_ (.I(_05846_),
    .Z(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11747_ (.I(_05768_),
    .Z(_05847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11748_ (.A1(_04223_),
    .A2(_05847_),
    .ZN(_05848_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11749_ (.I(_05848_),
    .Z(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11750_ (.I0(_05825_),
    .I1(\u2.mem[184][0] ),
    .S(_05849_),
    .Z(_05850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11751_ (.I(_05850_),
    .Z(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11752_ (.I0(_05829_),
    .I1(\u2.mem[184][1] ),
    .S(_05849_),
    .Z(_05851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11753_ (.I(_05851_),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11754_ (.I0(_05831_),
    .I1(\u2.mem[184][2] ),
    .S(_05849_),
    .Z(_05852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11755_ (.I(_05852_),
    .Z(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11756_ (.I0(_05833_),
    .I1(\u2.mem[184][3] ),
    .S(_05849_),
    .Z(_05853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11757_ (.I(_05853_),
    .Z(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11758_ (.I0(_05835_),
    .I1(\u2.mem[184][4] ),
    .S(_05848_),
    .Z(_05854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11759_ (.I(_05854_),
    .Z(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11760_ (.I0(_05837_),
    .I1(\u2.mem[184][5] ),
    .S(_05848_),
    .Z(_05855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11761_ (.I(_05855_),
    .Z(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11762_ (.A1(_04248_),
    .A2(_05847_),
    .ZN(_05856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11763_ (.I(_05856_),
    .Z(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11764_ (.I0(_05825_),
    .I1(\u2.mem[185][0] ),
    .S(_05857_),
    .Z(_05858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11765_ (.I(_05858_),
    .Z(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11766_ (.I0(_05829_),
    .I1(\u2.mem[185][1] ),
    .S(_05857_),
    .Z(_05859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11767_ (.I(_05859_),
    .Z(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11768_ (.I0(_05831_),
    .I1(\u2.mem[185][2] ),
    .S(_05857_),
    .Z(_05860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11769_ (.I(_05860_),
    .Z(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11770_ (.I0(_05833_),
    .I1(\u2.mem[185][3] ),
    .S(_05857_),
    .Z(_05861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11771_ (.I(_05861_),
    .Z(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11772_ (.I0(_05835_),
    .I1(\u2.mem[185][4] ),
    .S(_05856_),
    .Z(_05862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11773_ (.I(_05862_),
    .Z(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11774_ (.I0(_05837_),
    .I1(\u2.mem[185][5] ),
    .S(_05856_),
    .Z(_05863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11775_ (.I(_05863_),
    .Z(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11776_ (.I(_03655_),
    .Z(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11777_ (.A1(_04287_),
    .A2(_05847_),
    .ZN(_05865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11778_ (.I(_05865_),
    .Z(_05866_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11779_ (.I0(_05864_),
    .I1(\u2.mem[186][0] ),
    .S(_05866_),
    .Z(_05867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11780_ (.I(_05867_),
    .Z(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11781_ (.I(_03662_),
    .Z(_05868_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11782_ (.I0(_05868_),
    .I1(\u2.mem[186][1] ),
    .S(_05866_),
    .Z(_05869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11783_ (.I(_05869_),
    .Z(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11784_ (.I(_03666_),
    .Z(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11785_ (.I0(_05870_),
    .I1(\u2.mem[186][2] ),
    .S(_05866_),
    .Z(_05871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11786_ (.I(_05871_),
    .Z(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11787_ (.I(_03670_),
    .Z(_05872_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11788_ (.I0(_05872_),
    .I1(\u2.mem[186][3] ),
    .S(_05866_),
    .Z(_05873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11789_ (.I(_05873_),
    .Z(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11790_ (.I(_03674_),
    .Z(_05874_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11791_ (.I0(_05874_),
    .I1(\u2.mem[186][4] ),
    .S(_05865_),
    .Z(_05875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11792_ (.I(_05875_),
    .Z(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11793_ (.I(_03679_),
    .Z(_05876_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11794_ (.I0(_05876_),
    .I1(\u2.mem[186][5] ),
    .S(_05865_),
    .Z(_05877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11795_ (.I(_05877_),
    .Z(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11796_ (.A1(_04310_),
    .A2(_05847_),
    .ZN(_05878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11797_ (.I(_05878_),
    .Z(_05879_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11798_ (.I0(_05864_),
    .I1(\u2.mem[187][0] ),
    .S(_05879_),
    .Z(_05880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11799_ (.I(_05880_),
    .Z(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11800_ (.I0(_05868_),
    .I1(\u2.mem[187][1] ),
    .S(_05879_),
    .Z(_05881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11801_ (.I(_05881_),
    .Z(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11802_ (.I0(_05870_),
    .I1(\u2.mem[187][2] ),
    .S(_05879_),
    .Z(_05882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11803_ (.I(_05882_),
    .Z(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11804_ (.I0(_05872_),
    .I1(\u2.mem[187][3] ),
    .S(_05879_),
    .Z(_05883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11805_ (.I(_05883_),
    .Z(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11806_ (.I0(_05874_),
    .I1(\u2.mem[187][4] ),
    .S(_05878_),
    .Z(_05884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11807_ (.I(_05884_),
    .Z(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11808_ (.I0(_05876_),
    .I1(\u2.mem[187][5] ),
    .S(_05878_),
    .Z(_05885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11809_ (.I(_05885_),
    .Z(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11810_ (.I(_05768_),
    .Z(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11811_ (.A1(_04333_),
    .A2(_05886_),
    .ZN(_05887_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11812_ (.I(_05887_),
    .Z(_05888_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11813_ (.I0(_05864_),
    .I1(\u2.mem[188][0] ),
    .S(_05888_),
    .Z(_05889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11814_ (.I(_05889_),
    .Z(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11815_ (.I0(_05868_),
    .I1(\u2.mem[188][1] ),
    .S(_05888_),
    .Z(_05890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11816_ (.I(_05890_),
    .Z(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11817_ (.I0(_05870_),
    .I1(\u2.mem[188][2] ),
    .S(_05888_),
    .Z(_05891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11818_ (.I(_05891_),
    .Z(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11819_ (.I0(_05872_),
    .I1(\u2.mem[188][3] ),
    .S(_05888_),
    .Z(_05892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11820_ (.I(_05892_),
    .Z(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11821_ (.I0(_05874_),
    .I1(\u2.mem[188][4] ),
    .S(_05887_),
    .Z(_05893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11822_ (.I(_05893_),
    .Z(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11823_ (.I0(_05876_),
    .I1(\u2.mem[188][5] ),
    .S(_05887_),
    .Z(_05894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11824_ (.I(_05894_),
    .Z(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11825_ (.A1(_05411_),
    .A2(_05886_),
    .ZN(_05895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11826_ (.I(_05895_),
    .Z(_05896_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11827_ (.I0(_05864_),
    .I1(\u2.mem[189][0] ),
    .S(_05896_),
    .Z(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11828_ (.I(_05897_),
    .Z(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11829_ (.I0(_05868_),
    .I1(\u2.mem[189][1] ),
    .S(_05896_),
    .Z(_05898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11830_ (.I(_05898_),
    .Z(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11831_ (.I0(_05870_),
    .I1(\u2.mem[189][2] ),
    .S(_05896_),
    .Z(_05899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11832_ (.I(_05899_),
    .Z(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11833_ (.I0(_05872_),
    .I1(\u2.mem[189][3] ),
    .S(_05896_),
    .Z(_05900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11834_ (.I(_05900_),
    .Z(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11835_ (.I0(_05874_),
    .I1(\u2.mem[189][4] ),
    .S(_05895_),
    .Z(_05901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11836_ (.I(_05901_),
    .Z(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11837_ (.I0(_05876_),
    .I1(\u2.mem[189][5] ),
    .S(_05895_),
    .Z(_05902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11838_ (.I(_05902_),
    .Z(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11839_ (.I(_03655_),
    .Z(_05903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11840_ (.A1(_04393_),
    .A2(_05886_),
    .ZN(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11841_ (.I(_05904_),
    .Z(_05905_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11842_ (.I0(_05903_),
    .I1(\u2.mem[190][0] ),
    .S(_05905_),
    .Z(_05906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11843_ (.I(_05906_),
    .Z(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11844_ (.I(_03662_),
    .Z(_05907_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11845_ (.I0(_05907_),
    .I1(\u2.mem[190][1] ),
    .S(_05905_),
    .Z(_05908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11846_ (.I(_05908_),
    .Z(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11847_ (.I(_03666_),
    .Z(_05909_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11848_ (.I0(_05909_),
    .I1(\u2.mem[190][2] ),
    .S(_05905_),
    .Z(_05910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11849_ (.I(_05910_),
    .Z(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11850_ (.I(_03670_),
    .Z(_05911_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11851_ (.I0(_05911_),
    .I1(\u2.mem[190][3] ),
    .S(_05905_),
    .Z(_05912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11852_ (.I(_05912_),
    .Z(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11853_ (.I(_03674_),
    .Z(_05913_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11854_ (.I0(_05913_),
    .I1(\u2.mem[190][4] ),
    .S(_05904_),
    .Z(_05914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11855_ (.I(_05914_),
    .Z(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11856_ (.I(_03679_),
    .Z(_05915_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11857_ (.I0(_05915_),
    .I1(\u2.mem[190][5] ),
    .S(_05904_),
    .Z(_05916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11858_ (.I(_05916_),
    .Z(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11859_ (.A1(_04416_),
    .A2(_05886_),
    .ZN(_05917_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11860_ (.I(_05917_),
    .Z(_05918_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11861_ (.I0(_05903_),
    .I1(\u2.mem[191][0] ),
    .S(_05918_),
    .Z(_05919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11862_ (.I(_05919_),
    .Z(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11863_ (.I0(_05907_),
    .I1(\u2.mem[191][1] ),
    .S(_05918_),
    .Z(_05920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11864_ (.I(_05920_),
    .Z(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11865_ (.I0(_05909_),
    .I1(\u2.mem[191][2] ),
    .S(_05918_),
    .Z(_05921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11866_ (.I(_05921_),
    .Z(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11867_ (.I0(_05911_),
    .I1(\u2.mem[191][3] ),
    .S(_05918_),
    .Z(_05922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11868_ (.I(_05922_),
    .Z(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11869_ (.I0(_05913_),
    .I1(\u2.mem[191][4] ),
    .S(_05917_),
    .Z(_05923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11870_ (.I(_05923_),
    .Z(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11871_ (.I0(_05915_),
    .I1(\u2.mem[191][5] ),
    .S(_05917_),
    .Z(_05924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11872_ (.I(_05924_),
    .Z(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11873_ (.A1(\mem_address_trans[6].data_sync ),
    .A2(\mem_address_trans[7].data_sync ),
    .ZN(_05925_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11874_ (.A1(_03477_),
    .A2(\mem_address_trans[5].data_sync ),
    .A3(_05925_),
    .ZN(_05926_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11875_ (.A1(_03486_),
    .A2(_05926_),
    .Z(_05927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11876_ (.I(_05927_),
    .Z(_05928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11877_ (.I(_05928_),
    .Z(_05929_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11878_ (.I0(\u2.mem[192][0] ),
    .I1(_03492_),
    .S(_05929_),
    .Z(_05930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11879_ (.I(_05930_),
    .Z(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11880_ (.I0(\u2.mem[192][1] ),
    .I1(_03497_),
    .S(_05929_),
    .Z(_05931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11881_ (.I(_05931_),
    .Z(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11882_ (.I(_05928_),
    .Z(_05932_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11883_ (.I0(\u2.mem[192][2] ),
    .I1(_03500_),
    .S(_05932_),
    .Z(_05933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11884_ (.I(_05933_),
    .Z(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11885_ (.I0(\u2.mem[192][3] ),
    .I1(_03503_),
    .S(_05932_),
    .Z(_05934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11886_ (.I(_05934_),
    .Z(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11887_ (.I0(\u2.mem[192][4] ),
    .I1(_03507_),
    .S(_05932_),
    .Z(_05935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11888_ (.I(_05935_),
    .Z(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11889_ (.I0(\u2.mem[192][5] ),
    .I1(_03511_),
    .S(_05932_),
    .Z(_05936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11890_ (.I(_05936_),
    .Z(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11891_ (.I(_05928_),
    .Z(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11892_ (.I0(\u2.mem[192][6] ),
    .I1(_03513_),
    .S(_05937_),
    .Z(_05938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11893_ (.I(_05938_),
    .Z(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11894_ (.I0(\u2.mem[192][7] ),
    .I1(_03515_),
    .S(_05937_),
    .Z(_05939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11895_ (.I(_05939_),
    .Z(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11896_ (.I0(\u2.mem[192][8] ),
    .I1(_03518_),
    .S(_05937_),
    .Z(_05940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11897_ (.I(_05940_),
    .Z(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11898_ (.I0(\u2.mem[192][9] ),
    .I1(_03521_),
    .S(_05937_),
    .Z(_05941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11899_ (.I(_05941_),
    .Z(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11900_ (.I(_05927_),
    .Z(_05942_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11901_ (.I0(\u2.mem[192][10] ),
    .I1(_03523_),
    .S(_05942_),
    .Z(_05943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11902_ (.I(_05943_),
    .Z(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11903_ (.I0(\u2.mem[192][11] ),
    .I1(_03525_),
    .S(_05942_),
    .Z(_05944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11904_ (.I(_05944_),
    .Z(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11905_ (.I0(\u2.mem[192][12] ),
    .I1(_03528_),
    .S(_05942_),
    .Z(_05945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11906_ (.I(_05945_),
    .Z(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11907_ (.I0(\u2.mem[192][13] ),
    .I1(_03531_),
    .S(_05942_),
    .Z(_05946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11908_ (.I(_05946_),
    .Z(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11909_ (.I0(\u2.mem[192][14] ),
    .I1(_03533_),
    .S(_05928_),
    .Z(_05947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11910_ (.I(_05947_),
    .Z(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11911_ (.A1(_03535_),
    .A2(_05929_),
    .ZN(_05948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11912_ (.A1(_01981_),
    .A2(_05929_),
    .B(_05948_),
    .ZN(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11913_ (.A1(_04013_),
    .A2(_05926_),
    .ZN(_05949_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11914_ (.I(_05949_),
    .Z(_05950_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11915_ (.I0(_05903_),
    .I1(\u2.mem[193][0] ),
    .S(_05950_),
    .Z(_05951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11916_ (.I(_05951_),
    .Z(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11917_ (.I0(_05907_),
    .I1(\u2.mem[193][1] ),
    .S(_05950_),
    .Z(_05952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11918_ (.I(_05952_),
    .Z(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11919_ (.I0(_05909_),
    .I1(\u2.mem[193][2] ),
    .S(_05950_),
    .Z(_05953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11920_ (.I(_05953_),
    .Z(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11921_ (.I0(_05911_),
    .I1(\u2.mem[193][3] ),
    .S(_05950_),
    .Z(_05954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11922_ (.I(_05954_),
    .Z(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11923_ (.I(_05949_),
    .Z(_05955_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11924_ (.I0(_05913_),
    .I1(\u2.mem[193][4] ),
    .S(_05955_),
    .Z(_05956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11925_ (.I(_05956_),
    .Z(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11926_ (.I0(_05915_),
    .I1(\u2.mem[193][5] ),
    .S(_05955_),
    .Z(_05957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11927_ (.I(_05957_),
    .Z(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11928_ (.I0(_05209_),
    .I1(\u2.mem[193][6] ),
    .S(_05955_),
    .Z(_05958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11929_ (.I(_05958_),
    .Z(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11930_ (.I0(_05211_),
    .I1(\u2.mem[193][7] ),
    .S(_05955_),
    .Z(_05959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11931_ (.I(_05959_),
    .Z(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11932_ (.I(_05949_),
    .Z(_05960_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11933_ (.I0(_05213_),
    .I1(\u2.mem[193][8] ),
    .S(_05960_),
    .Z(_05961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11934_ (.I(_05961_),
    .Z(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11935_ (.I0(_05216_),
    .I1(\u2.mem[193][9] ),
    .S(_05960_),
    .Z(_05962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11936_ (.I(_05962_),
    .Z(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11937_ (.I0(_05218_),
    .I1(\u2.mem[193][10] ),
    .S(_05960_),
    .Z(_05963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11938_ (.I(_05963_),
    .Z(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11939_ (.I0(_05220_),
    .I1(\u2.mem[193][11] ),
    .S(_05960_),
    .Z(_05964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11940_ (.I(_05964_),
    .Z(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11941_ (.I(_05949_),
    .Z(_05965_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11942_ (.I0(_05222_),
    .I1(\u2.mem[193][12] ),
    .S(_05965_),
    .Z(_05966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11943_ (.I(_05966_),
    .Z(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11944_ (.I0(_05225_),
    .I1(\u2.mem[193][13] ),
    .S(_05965_),
    .Z(_05967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11945_ (.I(_05967_),
    .Z(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11946_ (.I0(_05227_),
    .I1(\u2.mem[193][14] ),
    .S(_05965_),
    .Z(_05968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11947_ (.I(_05968_),
    .Z(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11948_ (.I0(_05229_),
    .I1(\u2.mem[193][15] ),
    .S(_05965_),
    .Z(_05969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11949_ (.I(_05969_),
    .Z(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11950_ (.A1(_03582_),
    .A2(_05926_),
    .ZN(_05970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11951_ (.I(_05970_),
    .Z(_05971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11952_ (.I(_05971_),
    .Z(_05972_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11953_ (.I0(_05903_),
    .I1(\u2.mem[194][0] ),
    .S(_05972_),
    .Z(_05973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11954_ (.I(_05973_),
    .Z(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11955_ (.I0(_05907_),
    .I1(\u2.mem[194][1] ),
    .S(_05972_),
    .Z(_05974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11956_ (.I(_05974_),
    .Z(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11957_ (.I(_05971_),
    .Z(_05975_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11958_ (.I0(_05909_),
    .I1(\u2.mem[194][2] ),
    .S(_05975_),
    .Z(_05976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11959_ (.I(_05976_),
    .Z(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11960_ (.I0(_05911_),
    .I1(\u2.mem[194][3] ),
    .S(_05975_),
    .Z(_05977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11961_ (.I(_05977_),
    .Z(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11962_ (.I0(_05913_),
    .I1(\u2.mem[194][4] ),
    .S(_05975_),
    .Z(_05978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11963_ (.I(_05978_),
    .Z(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11964_ (.I0(_05915_),
    .I1(\u2.mem[194][5] ),
    .S(_05975_),
    .Z(_05979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11965_ (.I(_05979_),
    .Z(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11966_ (.I(_05971_),
    .Z(_05980_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11967_ (.I0(_05209_),
    .I1(\u2.mem[194][6] ),
    .S(_05980_),
    .Z(_05981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11968_ (.I(_05981_),
    .Z(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11969_ (.I0(_05211_),
    .I1(\u2.mem[194][7] ),
    .S(_05980_),
    .Z(_05982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11970_ (.I(_05982_),
    .Z(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11971_ (.I0(_05213_),
    .I1(\u2.mem[194][8] ),
    .S(_05980_),
    .Z(_05983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11972_ (.I(_05983_),
    .Z(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11973_ (.I0(_05216_),
    .I1(\u2.mem[194][9] ),
    .S(_05980_),
    .Z(_05984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11974_ (.I(_05984_),
    .Z(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11975_ (.I(_05970_),
    .Z(_05985_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11976_ (.I0(_05218_),
    .I1(\u2.mem[194][10] ),
    .S(_05985_),
    .Z(_05986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11977_ (.I(_05986_),
    .Z(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11978_ (.I0(_05220_),
    .I1(\u2.mem[194][11] ),
    .S(_05985_),
    .Z(_05987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11979_ (.I(_05987_),
    .Z(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11980_ (.I0(_05222_),
    .I1(\u2.mem[194][12] ),
    .S(_05985_),
    .Z(_05988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11981_ (.I(_05988_),
    .Z(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11982_ (.I0(_05225_),
    .I1(\u2.mem[194][13] ),
    .S(_05985_),
    .Z(_05989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11983_ (.I(_05989_),
    .Z(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11984_ (.I0(_05227_),
    .I1(\u2.mem[194][14] ),
    .S(_05971_),
    .Z(_05990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11985_ (.I(_05990_),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11986_ (.A1(_03535_),
    .A2(_05972_),
    .ZN(_05991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11987_ (.A1(_01979_),
    .A2(_05972_),
    .B(_05991_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11988_ (.D(_00000_),
    .CLK(clknet_leaf_362_clock),
    .Q(\u3.data ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11989_ (.D(_00001_),
    .CLK(clknet_leaf_318_clock),
    .Q(\u2.mem[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11990_ (.D(_00002_),
    .CLK(clknet_leaf_329_clock),
    .Q(\u2.mem[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11991_ (.D(_00003_),
    .CLK(clknet_leaf_318_clock),
    .Q(\u2.mem[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11992_ (.D(_00004_),
    .CLK(clknet_leaf_329_clock),
    .Q(\u2.mem[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11993_ (.D(_00005_),
    .CLK(clknet_leaf_318_clock),
    .Q(\u2.mem[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11994_ (.D(_00006_),
    .CLK(clknet_leaf_320_clock),
    .Q(\u2.mem[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11995_ (.D(_00007_),
    .CLK(clknet_leaf_319_clock),
    .Q(\u2.mem[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11996_ (.D(_00008_),
    .CLK(clknet_leaf_320_clock),
    .Q(\u2.mem[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11997_ (.D(_00009_),
    .CLK(clknet_leaf_33_clock),
    .Q(\u2.mem[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11998_ (.D(_00010_),
    .CLK(clknet_leaf_28_clock),
    .Q(\u2.mem[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11999_ (.D(_00011_),
    .CLK(clknet_leaf_28_clock),
    .Q(\u2.mem[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12000_ (.D(_00012_),
    .CLK(clknet_leaf_28_clock),
    .Q(\u2.mem[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12001_ (.D(_00013_),
    .CLK(clknet_leaf_42_clock),
    .Q(\u2.mem[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12002_ (.D(_00014_),
    .CLK(clknet_leaf_42_clock),
    .Q(\u2.mem[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12003_ (.D(_00015_),
    .CLK(clknet_leaf_41_clock),
    .Q(\u2.mem[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12004_ (.D(_00016_),
    .CLK(clknet_leaf_40_clock),
    .Q(\u2.mem[0][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12005_ (.D(net24),
    .CLK(clknet_2_3__leaf_clock_a),
    .Q(\mem_address_trans[0].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12006_ (.D(\mem_address_trans[0].A ),
    .CLK(clknet_leaf_312_clock),
    .Q(\mem_address_trans[0].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12007_ (.D(net25),
    .CLK(clknet_2_2__leaf_clock_a),
    .Q(\mem_address_trans[1].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12008_ (.D(\mem_address_trans[1].A ),
    .CLK(clknet_leaf_299_clock),
    .Q(\mem_address_trans[1].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12009_ (.D(net26),
    .CLK(clknet_2_0__leaf_clock_a),
    .Q(\mem_address_trans[2].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12010_ (.D(\mem_address_trans[2].A ),
    .CLK(clknet_leaf_312_clock),
    .Q(\mem_address_trans[2].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12011_ (.D(net27),
    .CLK(clknet_2_1__leaf_clock_a),
    .Q(\mem_address_trans[3].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12012_ (.D(\mem_address_trans[3].A ),
    .CLK(clknet_leaf_244_clock),
    .Q(\mem_address_trans[3].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12013_ (.D(net28),
    .CLK(clknet_2_0__leaf_clock_a),
    .Q(\mem_address_trans[4].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12014_ (.D(\mem_address_trans[4].A ),
    .CLK(clknet_leaf_289_clock),
    .Q(\mem_address_trans[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12015_ (.D(net29),
    .CLK(clknet_2_2__leaf_clock_a),
    .Q(\mem_address_trans[5].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12016_ (.D(\mem_address_trans[5].A ),
    .CLK(clknet_leaf_294_clock),
    .Q(\mem_address_trans[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12017_ (.D(net30),
    .CLK(clknet_2_2__leaf_clock_a),
    .Q(\mem_address_trans[6].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12018_ (.D(\mem_address_trans[6].A ),
    .CLK(clknet_leaf_299_clock),
    .Q(\mem_address_trans[6].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12019_ (.D(net31),
    .CLK(clknet_2_2__leaf_clock_a),
    .Q(\mem_address_trans[7].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12020_ (.D(\mem_address_trans[7].A ),
    .CLK(clknet_leaf_289_clock),
    .Q(\mem_address_trans[7].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12021_ (.D(net32),
    .CLK(clknet_2_1__leaf_clock_a),
    .Q(\mem_address_trans[8].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12022_ (.D(\mem_address_trans[8].A ),
    .CLK(clknet_leaf_287_clock),
    .Q(\mem_address_trans[8].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12023_ (.D(net33),
    .CLK(clknet_2_1__leaf_clock_a),
    .Q(\mem_address_trans[9].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12024_ (.D(\mem_address_trans[9].A ),
    .CLK(clknet_leaf_289_clock),
    .Q(\mem_address_trans[9].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12025_ (.D(net37),
    .CLK(clknet_2_3__leaf_clock_a),
    .Q(\row_select_trans[0].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12026_ (.D(\row_select_trans[0].A ),
    .CLK(clknet_leaf_302_clock),
    .Q(\row_select_trans[0].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12027_ (.D(net38),
    .CLK(clknet_2_0__leaf_clock_a),
    .Q(\row_select_trans[1].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12028_ (.D(\row_select_trans[1].A ),
    .CLK(clknet_leaf_307_clock),
    .Q(\row_select_trans[1].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12029_ (.D(net39),
    .CLK(clknet_2_2__leaf_clock_a),
    .Q(\row_select_trans[2].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12030_ (.D(\row_select_trans[2].A ),
    .CLK(clknet_leaf_307_clock),
    .Q(\row_select_trans[2].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12031_ (.D(net40),
    .CLK(clknet_2_3__leaf_clock_a),
    .Q(\row_select_trans[3].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12032_ (.D(\row_select_trans[3].A ),
    .CLK(clknet_leaf_302_clock),
    .Q(\row_select_trans[3].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12033_ (.D(net41),
    .CLK(clknet_2_3__leaf_clock_a),
    .Q(\row_select_trans[4].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12034_ (.D(\row_select_trans[4].A ),
    .CLK(clknet_leaf_289_clock),
    .Q(\row_select_trans[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12035_ (.D(net42),
    .CLK(clknet_2_3__leaf_clock_a),
    .Q(\row_select_trans[5].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12036_ (.D(\row_select_trans[5].A ),
    .CLK(clknet_leaf_311_clock),
    .Q(\row_select_trans[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12037_ (.D(net1),
    .CLK(clknet_2_0__leaf_clock_a),
    .Q(\col_select_trans[0].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12038_ (.D(\col_select_trans[0].A ),
    .CLK(clknet_leaf_302_clock),
    .Q(\col_select_trans[0].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12039_ (.D(net2),
    .CLK(clknet_2_2__leaf_clock_a),
    .Q(\col_select_trans[1].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12040_ (.D(\col_select_trans[1].A ),
    .CLK(clknet_leaf_299_clock),
    .Q(\col_select_trans[1].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12041_ (.D(net3),
    .CLK(clknet_2_3__leaf_clock_a),
    .Q(\col_select_trans[2].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12042_ (.D(\col_select_trans[2].A ),
    .CLK(clknet_leaf_299_clock),
    .Q(\col_select_trans[2].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12043_ (.D(net4),
    .CLK(clknet_2_2__leaf_clock_a),
    .Q(\col_select_trans[3].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12044_ (.D(\col_select_trans[3].A ),
    .CLK(clknet_leaf_299_clock),
    .Q(\col_select_trans[3].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12045_ (.D(net5),
    .CLK(clknet_2_2__leaf_clock_a),
    .Q(\col_select_trans[4].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12046_ (.D(\col_select_trans[4].A ),
    .CLK(clknet_leaf_288_clock),
    .Q(\col_select_trans[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12047_ (.D(net6),
    .CLK(clknet_2_2__leaf_clock_a),
    .Q(\col_select_trans[5].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12048_ (.D(\col_select_trans[5].A ),
    .CLK(clknet_leaf_288_clock),
    .Q(\col_select_trans[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12049_ (.D(net7),
    .CLK(clknet_2_3__leaf_clock_a),
    .Q(\data_in_trans[0].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12050_ (.D(\data_in_trans[0].A ),
    .CLK(clknet_leaf_288_clock),
    .Q(\data_in_trans[0].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12051_ (.D(net14),
    .CLK(clknet_2_0__leaf_clock_a),
    .Q(\data_in_trans[1].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12052_ (.D(\data_in_trans[1].A ),
    .CLK(clknet_leaf_287_clock),
    .Q(\data_in_trans[1].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12053_ (.D(net15),
    .CLK(clknet_2_0__leaf_clock_a),
    .Q(\data_in_trans[2].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12054_ (.D(\data_in_trans[2].A ),
    .CLK(clknet_leaf_287_clock),
    .Q(\data_in_trans[2].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12055_ (.D(net16),
    .CLK(clknet_2_2__leaf_clock_a),
    .Q(\data_in_trans[3].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12056_ (.D(\data_in_trans[3].A ),
    .CLK(clknet_leaf_288_clock),
    .Q(\data_in_trans[3].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12057_ (.D(net17),
    .CLK(clknet_2_1__leaf_clock_a),
    .Q(\data_in_trans[4].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12058_ (.D(\data_in_trans[4].A ),
    .CLK(clknet_leaf_300_clock),
    .Q(\data_in_trans[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12059_ (.D(net18),
    .CLK(clknet_2_1__leaf_clock_a),
    .Q(\data_in_trans[5].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12060_ (.D(\data_in_trans[5].A ),
    .CLK(clknet_leaf_300_clock),
    .Q(\data_in_trans[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12061_ (.D(net19),
    .CLK(clknet_2_0__leaf_clock_a),
    .Q(\data_in_trans[6].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12062_ (.D(\data_in_trans[6].A ),
    .CLK(clknet_leaf_302_clock),
    .Q(\data_in_trans[6].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12063_ (.D(net20),
    .CLK(clknet_2_3__leaf_clock_a),
    .Q(\data_in_trans[7].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12064_ (.D(\data_in_trans[7].A ),
    .CLK(clknet_leaf_300_clock),
    .Q(\data_in_trans[7].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12065_ (.D(net21),
    .CLK(clknet_2_3__leaf_clock_a),
    .Q(\data_in_trans[8].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12066_ (.D(\data_in_trans[8].A ),
    .CLK(clknet_leaf_32_clock),
    .Q(\data_in_trans[8].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12067_ (.D(net22),
    .CLK(clknet_2_1__leaf_clock_a),
    .Q(\data_in_trans[9].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12068_ (.D(\data_in_trans[9].A ),
    .CLK(clknet_leaf_33_clock),
    .Q(\data_in_trans[9].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12069_ (.D(net8),
    .CLK(clknet_2_0__leaf_clock_a),
    .Q(\data_in_trans[10].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12070_ (.D(\data_in_trans[10].A ),
    .CLK(clknet_leaf_28_clock),
    .Q(\data_in_trans[10].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12071_ (.D(net9),
    .CLK(clknet_2_1__leaf_clock_a),
    .Q(\data_in_trans[11].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12072_ (.D(\data_in_trans[11].A ),
    .CLK(clknet_leaf_28_clock),
    .Q(\data_in_trans[11].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12073_ (.D(net10),
    .CLK(clknet_2_1__leaf_clock_a),
    .Q(\data_in_trans[12].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12074_ (.D(\data_in_trans[12].A ),
    .CLK(clknet_leaf_343_clock),
    .Q(\data_in_trans[12].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12075_ (.D(net11),
    .CLK(clknet_2_2__leaf_clock_a),
    .Q(\data_in_trans[13].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12076_ (.D(\data_in_trans[13].A ),
    .CLK(clknet_leaf_343_clock),
    .Q(\data_in_trans[13].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12077_ (.D(net12),
    .CLK(clknet_2_2__leaf_clock_a),
    .Q(\data_in_trans[14].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12078_ (.D(\data_in_trans[14].A ),
    .CLK(clknet_leaf_343_clock),
    .Q(\data_in_trans[14].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12079_ (.D(net13),
    .CLK(clknet_2_1__leaf_clock_a),
    .Q(\data_in_trans[15].A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12080_ (.D(\data_in_trans[15].A ),
    .CLK(clknet_leaf_303_clock),
    .Q(\data_in_trans[15].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12081_ (.D(net45),
    .CLK(clknet_leaf_362_clock),
    .Q(\output_active_hold[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12082_ (.D(\output_active_hold[0] ),
    .CLK(clknet_leaf_363_clock),
    .Q(\output_active_hold[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12083_ (.D(\output_active_hold[1] ),
    .CLK(clknet_leaf_363_clock),
    .Q(\output_active_hold[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12084_ (.D(\output_active_hold[2] ),
    .CLK(clknet_leaf_363_clock),
    .Q(\output_active_hold[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12085_ (.D(net34),
    .CLK(clknet_2_2__leaf_clock_a),
    .Q(\mem_write_n_trans.A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12086_ (.D(\mem_write_n_trans.A ),
    .CLK(clknet_leaf_288_clock),
    .Q(\mem_write_n_trans.data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12087_ (.D(net36),
    .CLK(clknet_2_1__leaf_clock_a),
    .Q(\row_col_select_trans.A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12088_ (.D(\row_col_select_trans.A ),
    .CLK(clknet_leaf_298_clock),
    .Q(\row_col_select_trans.data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12089_ (.D(net35),
    .CLK(clknet_2_0__leaf_clock_a),
    .Q(\output_active_trans.A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12090_ (.D(\output_active_trans.A ),
    .CLK(clknet_leaf_303_clock),
    .Q(\output_active_trans.data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12091_ (.D(net23),
    .CLK(clknet_2_3__leaf_clock_a),
    .Q(\inverter_select_trans.A ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12092_ (.D(\inverter_select_trans.A ),
    .CLK(clknet_leaf_302_clock),
    .Q(\inverter_select_trans.data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12093_ (.D(_00017_),
    .CLK(clknet_leaf_363_clock),
    .Q(\u3.enable ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12094_ (.D(_01486_),
    .CLK(clknet_leaf_218_clock),
    .Q(\u2.active_mem[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12095_ (.D(_01493_),
    .CLK(clknet_leaf_214_clock),
    .Q(\u2.active_mem[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12096_ (.D(_01494_),
    .CLK(clknet_leaf_214_clock),
    .Q(\u2.active_mem[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12097_ (.D(_01495_),
    .CLK(clknet_leaf_219_clock),
    .Q(\u2.active_mem[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12098_ (.D(_01496_),
    .CLK(clknet_leaf_224_clock),
    .Q(\u2.active_mem[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12099_ (.D(_01497_),
    .CLK(clknet_leaf_149_clock),
    .Q(\u2.active_mem[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12100_ (.D(_01498_),
    .CLK(clknet_leaf_149_clock),
    .Q(\u2.active_mem[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12101_ (.D(_01499_),
    .CLK(clknet_leaf_144_clock),
    .Q(\u2.active_mem[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12102_ (.D(_01500_),
    .CLK(clknet_leaf_62_clock),
    .Q(\u2.active_mem[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12103_ (.D(_01501_),
    .CLK(clknet_leaf_62_clock),
    .Q(\u2.active_mem[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12104_ (.D(_01487_),
    .CLK(clknet_leaf_63_clock),
    .Q(\u2.active_mem[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12105_ (.D(_01488_),
    .CLK(clknet_leaf_63_clock),
    .Q(\u2.active_mem[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12106_ (.D(_01489_),
    .CLK(clknet_leaf_58_clock),
    .Q(\u2.active_mem[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12107_ (.D(_01490_),
    .CLK(clknet_leaf_135_clock),
    .Q(\u2.active_mem[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12108_ (.D(_01491_),
    .CLK(clknet_leaf_135_clock),
    .Q(\u2.active_mem[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12109_ (.D(_01492_),
    .CLK(clknet_leaf_140_clock),
    .Q(\u2.active_mem[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12110_ (.D(_05992_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u2.driver_enable ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12111_ (.D(_01474_),
    .CLK(clknet_leaf_332_clock),
    .Q(\u2.select_mem_row[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12112_ (.D(_01475_),
    .CLK(clknet_leaf_334_clock),
    .Q(\u2.select_mem_row[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12113_ (.D(_01476_),
    .CLK(clknet_leaf_331_clock),
    .Q(\u2.select_mem_row[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12114_ (.D(_01477_),
    .CLK(clknet_leaf_333_clock),
    .Q(\u2.select_mem_row[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12115_ (.D(_01478_),
    .CLK(clknet_leaf_332_clock),
    .Q(\u2.select_mem_row[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12116_ (.D(_01479_),
    .CLK(clknet_leaf_328_clock),
    .Q(\u2.select_mem_row[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12117_ (.D(_01480_),
    .CLK(clknet_leaf_332_clock),
    .Q(\u2.select_mem_col[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12118_ (.D(_01481_),
    .CLK(clknet_leaf_334_clock),
    .Q(\u2.select_mem_col[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12119_ (.D(_01482_),
    .CLK(clknet_leaf_332_clock),
    .Q(\u2.select_mem_col[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12120_ (.D(_01483_),
    .CLK(clknet_leaf_333_clock),
    .Q(\u2.select_mem_col[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12121_ (.D(_01484_),
    .CLK(clknet_leaf_328_clock),
    .Q(\u2.select_mem_col[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12122_ (.D(_01485_),
    .CLK(clknet_leaf_328_clock),
    .Q(\u2.select_mem_col[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12123_ (.D(_01458_),
    .CLK(clknet_leaf_37_clock),
    .Q(\u2.driver_mem[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12124_ (.D(_01465_),
    .CLK(clknet_leaf_36_clock),
    .Q(\u2.driver_mem[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12125_ (.D(_01466_),
    .CLK(clknet_leaf_334_clock),
    .Q(\u2.driver_mem[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12126_ (.D(_01467_),
    .CLK(clknet_leaf_336_clock),
    .Q(\u2.driver_mem[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12127_ (.D(_01468_),
    .CLK(clknet_leaf_36_clock),
    .Q(\u2.driver_mem[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12128_ (.D(_01469_),
    .CLK(clknet_leaf_37_clock),
    .Q(\u2.driver_mem[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12129_ (.D(_01470_),
    .CLK(clknet_leaf_35_clock),
    .Q(\u2.driver_mem[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12130_ (.D(_01471_),
    .CLK(clknet_leaf_35_clock),
    .Q(\u2.driver_mem[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12131_ (.D(_01472_),
    .CLK(clknet_leaf_35_clock),
    .Q(\u2.driver_mem[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12132_ (.D(_01473_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u2.driver_mem[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12133_ (.D(_01459_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u2.driver_mem[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12134_ (.D(_01460_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u2.driver_mem[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12135_ (.D(_01461_),
    .CLK(clknet_leaf_37_clock),
    .Q(\u2.driver_mem[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12136_ (.D(_01462_),
    .CLK(clknet_leaf_37_clock),
    .Q(\u2.driver_mem[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12137_ (.D(_01463_),
    .CLK(clknet_leaf_38_clock),
    .Q(\u2.driver_mem[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12138_ (.D(_01464_),
    .CLK(clknet_leaf_38_clock),
    .Q(\u2.driver_mem[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12139_ (.D(_00018_),
    .CLK(clknet_leaf_212_clock),
    .Q(\u2.mem[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12140_ (.D(_00019_),
    .CLK(clknet_leaf_211_clock),
    .Q(\u2.mem[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12141_ (.D(_00020_),
    .CLK(clknet_leaf_211_clock),
    .Q(\u2.mem[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12142_ (.D(_00021_),
    .CLK(clknet_leaf_211_clock),
    .Q(\u2.mem[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12143_ (.D(_00022_),
    .CLK(clknet_leaf_218_clock),
    .Q(\u2.mem[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12144_ (.D(_00023_),
    .CLK(clknet_leaf_226_clock),
    .Q(\u2.mem[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12145_ (.D(_00024_),
    .CLK(clknet_leaf_218_clock),
    .Q(\u2.mem[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12146_ (.D(_00025_),
    .CLK(clknet_leaf_225_clock),
    .Q(\u2.mem[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12147_ (.D(_00026_),
    .CLK(clknet_leaf_73_clock),
    .Q(\u2.mem[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12148_ (.D(_00027_),
    .CLK(clknet_leaf_74_clock),
    .Q(\u2.mem[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12149_ (.D(_00028_),
    .CLK(clknet_leaf_73_clock),
    .Q(\u2.mem[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12150_ (.D(_00029_),
    .CLK(clknet_leaf_73_clock),
    .Q(\u2.mem[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12151_ (.D(_00030_),
    .CLK(clknet_leaf_64_clock),
    .Q(\u2.mem[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12152_ (.D(_00031_),
    .CLK(clknet_leaf_64_clock),
    .Q(\u2.mem[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12153_ (.D(_00032_),
    .CLK(clknet_leaf_56_clock),
    .Q(\u2.mem[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12154_ (.D(_00033_),
    .CLK(clknet_leaf_56_clock),
    .Q(\u2.mem[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12155_ (.D(_00034_),
    .CLK(clknet_leaf_204_clock),
    .Q(\u2.mem[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12156_ (.D(_00035_),
    .CLK(clknet_leaf_205_clock),
    .Q(\u2.mem[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12157_ (.D(_00036_),
    .CLK(clknet_leaf_205_clock),
    .Q(\u2.mem[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12158_ (.D(_00037_),
    .CLK(clknet_leaf_205_clock),
    .Q(\u2.mem[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12159_ (.D(_00038_),
    .CLK(clknet_leaf_153_clock),
    .Q(\u2.mem[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12160_ (.D(_00039_),
    .CLK(clknet_leaf_152_clock),
    .Q(\u2.mem[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12161_ (.D(_00040_),
    .CLK(clknet_leaf_154_clock),
    .Q(\u2.mem[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12162_ (.D(_00041_),
    .CLK(clknet_leaf_153_clock),
    .Q(\u2.mem[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12163_ (.D(_00042_),
    .CLK(clknet_leaf_91_clock),
    .Q(\u2.mem[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12164_ (.D(_00043_),
    .CLK(clknet_leaf_91_clock),
    .Q(\u2.mem[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12165_ (.D(_00044_),
    .CLK(clknet_leaf_91_clock),
    .Q(\u2.mem[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12166_ (.D(_00045_),
    .CLK(clknet_leaf_91_clock),
    .Q(\u2.mem[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12167_ (.D(_00046_),
    .CLK(clknet_leaf_109_clock),
    .Q(\u2.mem[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12168_ (.D(_00047_),
    .CLK(clknet_leaf_109_clock),
    .Q(\u2.mem[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12169_ (.D(_00048_),
    .CLK(clknet_leaf_131_clock),
    .Q(\u2.mem[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12170_ (.D(_00049_),
    .CLK(clknet_leaf_109_clock),
    .Q(\u2.mem[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12171_ (.D(_00050_),
    .CLK(clknet_leaf_209_clock),
    .Q(\u2.mem[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12172_ (.D(_00051_),
    .CLK(clknet_leaf_210_clock),
    .Q(\u2.mem[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12173_ (.D(_00052_),
    .CLK(clknet_leaf_210_clock),
    .Q(\u2.mem[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12174_ (.D(_00053_),
    .CLK(clknet_leaf_210_clock),
    .Q(\u2.mem[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12175_ (.D(_00054_),
    .CLK(clknet_leaf_218_clock),
    .Q(\u2.mem[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12176_ (.D(_00055_),
    .CLK(clknet_leaf_226_clock),
    .Q(\u2.mem[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12177_ (.D(_00056_),
    .CLK(clknet_leaf_218_clock),
    .Q(\u2.mem[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12178_ (.D(_00057_),
    .CLK(clknet_leaf_225_clock),
    .Q(\u2.mem[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12179_ (.D(_00058_),
    .CLK(clknet_leaf_76_clock),
    .Q(\u2.mem[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12180_ (.D(_00059_),
    .CLK(clknet_leaf_75_clock),
    .Q(\u2.mem[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12181_ (.D(_00060_),
    .CLK(clknet_leaf_77_clock),
    .Q(\u2.mem[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12182_ (.D(_00061_),
    .CLK(clknet_leaf_77_clock),
    .Q(\u2.mem[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12183_ (.D(_00062_),
    .CLK(clknet_leaf_61_clock),
    .Q(\u2.mem[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12184_ (.D(_00063_),
    .CLK(clknet_leaf_59_clock),
    .Q(\u2.mem[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12185_ (.D(_00064_),
    .CLK(clknet_leaf_59_clock),
    .Q(\u2.mem[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12186_ (.D(_00065_),
    .CLK(clknet_leaf_59_clock),
    .Q(\u2.mem[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12187_ (.D(_00066_),
    .CLK(clknet_leaf_251_clock),
    .Q(\u2.mem[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12188_ (.D(_00067_),
    .CLK(clknet_leaf_252_clock),
    .Q(\u2.mem[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12189_ (.D(_00068_),
    .CLK(clknet_leaf_252_clock),
    .Q(\u2.mem[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12190_ (.D(_00069_),
    .CLK(clknet_leaf_252_clock),
    .Q(\u2.mem[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12191_ (.D(_00070_),
    .CLK(clknet_leaf_237_clock),
    .Q(\u2.mem[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12192_ (.D(_00071_),
    .CLK(clknet_leaf_228_clock),
    .Q(\u2.mem[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12193_ (.D(_00072_),
    .CLK(clknet_leaf_228_clock),
    .Q(\u2.mem[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12194_ (.D(_00073_),
    .CLK(clknet_leaf_238_clock),
    .Q(\u2.mem[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12195_ (.D(_00074_),
    .CLK(clknet_leaf_72_clock),
    .Q(\u2.mem[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12196_ (.D(_00075_),
    .CLK(clknet_leaf_71_clock),
    .Q(\u2.mem[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12197_ (.D(_00076_),
    .CLK(clknet_leaf_72_clock),
    .Q(\u2.mem[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12198_ (.D(_00077_),
    .CLK(clknet_leaf_73_clock),
    .Q(\u2.mem[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12199_ (.D(_00078_),
    .CLK(clknet_leaf_66_clock),
    .Q(\u2.mem[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12200_ (.D(_00079_),
    .CLK(clknet_leaf_65_clock),
    .Q(\u2.mem[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12201_ (.D(_00080_),
    .CLK(clknet_leaf_54_clock),
    .Q(\u2.mem[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12202_ (.D(_00081_),
    .CLK(clknet_leaf_54_clock),
    .Q(\u2.mem[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12203_ (.D(_00082_),
    .CLK(clknet_leaf_217_clock),
    .Q(\u2.mem[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12204_ (.D(_00083_),
    .CLK(clknet_leaf_211_clock),
    .Q(\u2.mem[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12205_ (.D(_00084_),
    .CLK(clknet_leaf_212_clock),
    .Q(\u2.mem[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12206_ (.D(_00085_),
    .CLK(clknet_leaf_212_clock),
    .Q(\u2.mem[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12207_ (.D(_00086_),
    .CLK(clknet_leaf_229_clock),
    .Q(\u2.mem[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12208_ (.D(_00087_),
    .CLK(clknet_leaf_231_clock),
    .Q(\u2.mem[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12209_ (.D(_00088_),
    .CLK(clknet_leaf_232_clock),
    .Q(\u2.mem[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12210_ (.D(_00089_),
    .CLK(clknet_leaf_232_clock),
    .Q(\u2.mem[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12211_ (.D(_00090_),
    .CLK(clknet_leaf_65_clock),
    .Q(\u2.mem[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12212_ (.D(_00091_),
    .CLK(clknet_leaf_67_clock),
    .Q(\u2.mem[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12213_ (.D(_00092_),
    .CLK(clknet_leaf_68_clock),
    .Q(\u2.mem[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12214_ (.D(_00093_),
    .CLK(clknet_leaf_68_clock),
    .Q(\u2.mem[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12215_ (.D(_00094_),
    .CLK(clknet_leaf_53_clock),
    .Q(\u2.mem[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12216_ (.D(_00095_),
    .CLK(clknet_leaf_51_clock),
    .Q(\u2.mem[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12217_ (.D(_00096_),
    .CLK(clknet_leaf_53_clock),
    .Q(\u2.mem[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12218_ (.D(_00097_),
    .CLK(clknet_leaf_52_clock),
    .Q(\u2.mem[5][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12219_ (.D(_00098_),
    .CLK(clknet_leaf_217_clock),
    .Q(\u2.mem[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12220_ (.D(_00099_),
    .CLK(clknet_leaf_215_clock),
    .Q(\u2.mem[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12221_ (.D(_00100_),
    .CLK(clknet_leaf_213_clock),
    .Q(\u2.mem[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12222_ (.D(_00101_),
    .CLK(clknet_leaf_216_clock),
    .Q(\u2.mem[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12223_ (.D(_00102_),
    .CLK(clknet_leaf_231_clock),
    .Q(\u2.mem[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12224_ (.D(_00103_),
    .CLK(clknet_leaf_231_clock),
    .Q(\u2.mem[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12225_ (.D(_00104_),
    .CLK(clknet_leaf_232_clock),
    .Q(\u2.mem[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12226_ (.D(_00105_),
    .CLK(clknet_leaf_143_clock),
    .Q(\u2.mem[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12227_ (.D(_00106_),
    .CLK(clknet_leaf_64_clock),
    .Q(\u2.mem[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12228_ (.D(_00107_),
    .CLK(clknet_leaf_64_clock),
    .Q(\u2.mem[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12229_ (.D(_00108_),
    .CLK(clknet_leaf_69_clock),
    .Q(\u2.mem[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12230_ (.D(_00109_),
    .CLK(clknet_leaf_69_clock),
    .Q(\u2.mem[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12231_ (.D(_00110_),
    .CLK(clknet_leaf_52_clock),
    .Q(\u2.mem[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12232_ (.D(_00111_),
    .CLK(clknet_leaf_57_clock),
    .Q(\u2.mem[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12233_ (.D(_00112_),
    .CLK(clknet_leaf_57_clock),
    .Q(\u2.mem[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12234_ (.D(_00113_),
    .CLK(clknet_leaf_52_clock),
    .Q(\u2.mem[6][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12235_ (.D(_00114_),
    .CLK(clknet_leaf_211_clock),
    .Q(\u2.mem[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12236_ (.D(_00115_),
    .CLK(clknet_leaf_211_clock),
    .Q(\u2.mem[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12237_ (.D(_00116_),
    .CLK(clknet_leaf_211_clock),
    .Q(\u2.mem[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12238_ (.D(_00117_),
    .CLK(clknet_leaf_211_clock),
    .Q(\u2.mem[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12239_ (.D(_00118_),
    .CLK(clknet_leaf_217_clock),
    .Q(\u2.mem[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12240_ (.D(_00119_),
    .CLK(clknet_leaf_227_clock),
    .Q(\u2.mem[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12241_ (.D(_00120_),
    .CLK(clknet_leaf_227_clock),
    .Q(\u2.mem[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12242_ (.D(_00121_),
    .CLK(clknet_leaf_226_clock),
    .Q(\u2.mem[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12243_ (.D(_00122_),
    .CLK(clknet_leaf_73_clock),
    .Q(\u2.mem[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12244_ (.D(_00123_),
    .CLK(clknet_leaf_74_clock),
    .Q(\u2.mem[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12245_ (.D(_00124_),
    .CLK(clknet_leaf_73_clock),
    .Q(\u2.mem[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12246_ (.D(_00125_),
    .CLK(clknet_leaf_73_clock),
    .Q(\u2.mem[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12247_ (.D(_00126_),
    .CLK(clknet_leaf_55_clock),
    .Q(\u2.mem[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12248_ (.D(_00127_),
    .CLK(clknet_leaf_55_clock),
    .Q(\u2.mem[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12249_ (.D(_00128_),
    .CLK(clknet_leaf_55_clock),
    .Q(\u2.mem[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12250_ (.D(_00129_),
    .CLK(clknet_leaf_57_clock),
    .Q(\u2.mem[7][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12251_ (.D(_00130_),
    .CLK(clknet_leaf_216_clock),
    .Q(\u2.mem[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12252_ (.D(_00131_),
    .CLK(clknet_leaf_215_clock),
    .Q(\u2.mem[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12253_ (.D(_00132_),
    .CLK(clknet_leaf_213_clock),
    .Q(\u2.mem[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12254_ (.D(_00133_),
    .CLK(clknet_leaf_216_clock),
    .Q(\u2.mem[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12255_ (.D(_00134_),
    .CLK(clknet_leaf_217_clock),
    .Q(\u2.mem[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12256_ (.D(_00135_),
    .CLK(clknet_leaf_228_clock),
    .Q(\u2.mem[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12257_ (.D(_00136_),
    .CLK(clknet_leaf_228_clock),
    .Q(\u2.mem[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12258_ (.D(_00137_),
    .CLK(clknet_leaf_228_clock),
    .Q(\u2.mem[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12259_ (.D(_00138_),
    .CLK(clknet_leaf_70_clock),
    .Q(\u2.mem[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12260_ (.D(_00139_),
    .CLK(clknet_leaf_70_clock),
    .Q(\u2.mem[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12261_ (.D(_00140_),
    .CLK(clknet_leaf_70_clock),
    .Q(\u2.mem[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12262_ (.D(_00141_),
    .CLK(clknet_leaf_69_clock),
    .Q(\u2.mem[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12263_ (.D(_00142_),
    .CLK(clknet_leaf_55_clock),
    .Q(\u2.mem[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12264_ (.D(_00143_),
    .CLK(clknet_leaf_65_clock),
    .Q(\u2.mem[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12265_ (.D(_00144_),
    .CLK(clknet_leaf_54_clock),
    .Q(\u2.mem[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12266_ (.D(_00145_),
    .CLK(clknet_leaf_55_clock),
    .Q(\u2.mem[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12267_ (.D(_00146_),
    .CLK(clknet_leaf_184_clock),
    .Q(\u2.mem[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12268_ (.D(_00147_),
    .CLK(clknet_leaf_185_clock),
    .Q(\u2.mem[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12269_ (.D(_00148_),
    .CLK(clknet_leaf_185_clock),
    .Q(\u2.mem[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12270_ (.D(_00149_),
    .CLK(clknet_leaf_185_clock),
    .Q(\u2.mem[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12271_ (.D(_00150_),
    .CLK(clknet_leaf_166_clock),
    .Q(\u2.mem[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12272_ (.D(_00151_),
    .CLK(clknet_leaf_166_clock),
    .Q(\u2.mem[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12273_ (.D(_00152_),
    .CLK(clknet_leaf_165_clock),
    .Q(\u2.mem[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12274_ (.D(_00153_),
    .CLK(clknet_leaf_166_clock),
    .Q(\u2.mem[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12275_ (.D(_00154_),
    .CLK(clknet_leaf_102_clock),
    .Q(\u2.mem[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12276_ (.D(_00155_),
    .CLK(clknet_leaf_102_clock),
    .Q(\u2.mem[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12277_ (.D(_00156_),
    .CLK(clknet_leaf_102_clock),
    .Q(\u2.mem[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12278_ (.D(_00157_),
    .CLK(clknet_leaf_101_clock),
    .Q(\u2.mem[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12279_ (.D(_00158_),
    .CLK(clknet_leaf_120_clock),
    .Q(\u2.mem[9][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12280_ (.D(_00159_),
    .CLK(clknet_leaf_120_clock),
    .Q(\u2.mem[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12281_ (.D(_00160_),
    .CLK(clknet_leaf_119_clock),
    .Q(\u2.mem[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12282_ (.D(_00161_),
    .CLK(clknet_leaf_119_clock),
    .Q(\u2.mem[9][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12283_ (.D(_00162_),
    .CLK(clknet_leaf_184_clock),
    .Q(\u2.mem[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12284_ (.D(_00163_),
    .CLK(clknet_leaf_185_clock),
    .Q(\u2.mem[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12285_ (.D(_00164_),
    .CLK(clknet_leaf_185_clock),
    .Q(\u2.mem[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12286_ (.D(_00165_),
    .CLK(clknet_leaf_185_clock),
    .Q(\u2.mem[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12287_ (.D(_00166_),
    .CLK(clknet_leaf_164_clock),
    .Q(\u2.mem[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12288_ (.D(_00167_),
    .CLK(clknet_leaf_165_clock),
    .Q(\u2.mem[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12289_ (.D(_00168_),
    .CLK(clknet_leaf_165_clock),
    .Q(\u2.mem[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12290_ (.D(_00169_),
    .CLK(clknet_leaf_165_clock),
    .Q(\u2.mem[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12291_ (.D(_00170_),
    .CLK(clknet_leaf_103_clock),
    .Q(\u2.mem[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12292_ (.D(_00171_),
    .CLK(clknet_leaf_101_clock),
    .Q(\u2.mem[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12293_ (.D(_00172_),
    .CLK(clknet_leaf_101_clock),
    .Q(\u2.mem[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12294_ (.D(_00173_),
    .CLK(clknet_leaf_101_clock),
    .Q(\u2.mem[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12295_ (.D(_00174_),
    .CLK(clknet_leaf_120_clock),
    .Q(\u2.mem[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12296_ (.D(_00175_),
    .CLK(clknet_leaf_120_clock),
    .Q(\u2.mem[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12297_ (.D(_00176_),
    .CLK(clknet_leaf_120_clock),
    .Q(\u2.mem[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12298_ (.D(_00177_),
    .CLK(clknet_leaf_165_clock),
    .Q(\u2.mem[10][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12299_ (.D(_00178_),
    .CLK(clknet_leaf_170_clock),
    .Q(\u2.mem[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12300_ (.D(_00179_),
    .CLK(clknet_leaf_181_clock),
    .Q(\u2.mem[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12301_ (.D(_00180_),
    .CLK(clknet_leaf_183_clock),
    .Q(\u2.mem[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12302_ (.D(_00181_),
    .CLK(clknet_leaf_181_clock),
    .Q(\u2.mem[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12303_ (.D(_00182_),
    .CLK(clknet_leaf_166_clock),
    .Q(\u2.mem[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12304_ (.D(_00183_),
    .CLK(clknet_leaf_164_clock),
    .Q(\u2.mem[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12305_ (.D(_00184_),
    .CLK(clknet_leaf_164_clock),
    .Q(\u2.mem[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12306_ (.D(_00185_),
    .CLK(clknet_leaf_166_clock),
    .Q(\u2.mem[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12307_ (.D(_00186_),
    .CLK(clknet_leaf_104_clock),
    .Q(\u2.mem[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12308_ (.D(_00187_),
    .CLK(clknet_leaf_100_clock),
    .Q(\u2.mem[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12309_ (.D(_00188_),
    .CLK(clknet_leaf_100_clock),
    .Q(\u2.mem[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12310_ (.D(_00189_),
    .CLK(clknet_leaf_99_clock),
    .Q(\u2.mem[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12311_ (.D(_00190_),
    .CLK(clknet_leaf_118_clock),
    .Q(\u2.mem[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12312_ (.D(_00191_),
    .CLK(clknet_leaf_121_clock),
    .Q(\u2.mem[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12313_ (.D(_00192_),
    .CLK(clknet_leaf_118_clock),
    .Q(\u2.mem[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12314_ (.D(_00193_),
    .CLK(clknet_leaf_118_clock),
    .Q(\u2.mem[11][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12315_ (.D(_00194_),
    .CLK(clknet_leaf_222_clock),
    .Q(\u2.mem[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12316_ (.D(_00195_),
    .CLK(clknet_leaf_200_clock),
    .Q(\u2.mem[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12317_ (.D(_00196_),
    .CLK(clknet_leaf_197_clock),
    .Q(\u2.mem[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12318_ (.D(_00197_),
    .CLK(clknet_leaf_199_clock),
    .Q(\u2.mem[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12319_ (.D(_00198_),
    .CLK(clknet_leaf_157_clock),
    .Q(\u2.mem[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12320_ (.D(_00199_),
    .CLK(clknet_leaf_158_clock),
    .Q(\u2.mem[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12321_ (.D(_00200_),
    .CLK(clknet_leaf_158_clock),
    .Q(\u2.mem[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12322_ (.D(_00201_),
    .CLK(clknet_leaf_158_clock),
    .Q(\u2.mem[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12323_ (.D(_00202_),
    .CLK(clknet_leaf_84_clock),
    .Q(\u2.mem[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12324_ (.D(_00203_),
    .CLK(clknet_leaf_84_clock),
    .Q(\u2.mem[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12325_ (.D(_00204_),
    .CLK(clknet_leaf_85_clock),
    .Q(\u2.mem[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12326_ (.D(_00205_),
    .CLK(clknet_leaf_85_clock),
    .Q(\u2.mem[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12327_ (.D(_00206_),
    .CLK(clknet_leaf_126_clock),
    .Q(\u2.mem[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12328_ (.D(_00207_),
    .CLK(clknet_leaf_126_clock),
    .Q(\u2.mem[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12329_ (.D(_00208_),
    .CLK(clknet_leaf_125_clock),
    .Q(\u2.mem[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12330_ (.D(_00209_),
    .CLK(clknet_leaf_125_clock),
    .Q(\u2.mem[12][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12331_ (.D(_00210_),
    .CLK(clknet_leaf_207_clock),
    .Q(\u2.mem[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12332_ (.D(_00211_),
    .CLK(clknet_leaf_206_clock),
    .Q(\u2.mem[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12333_ (.D(_00212_),
    .CLK(clknet_leaf_209_clock),
    .Q(\u2.mem[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12334_ (.D(_00213_),
    .CLK(clknet_leaf_206_clock),
    .Q(\u2.mem[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12335_ (.D(_00214_),
    .CLK(clknet_leaf_152_clock),
    .Q(\u2.mem[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12336_ (.D(_00215_),
    .CLK(clknet_leaf_222_clock),
    .Q(\u2.mem[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12337_ (.D(_00216_),
    .CLK(clknet_leaf_152_clock),
    .Q(\u2.mem[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12338_ (.D(_00217_),
    .CLK(clknet_leaf_152_clock),
    .Q(\u2.mem[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12339_ (.D(_00218_),
    .CLK(clknet_leaf_77_clock),
    .Q(\u2.mem[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12340_ (.D(_00219_),
    .CLK(clknet_leaf_80_clock),
    .Q(\u2.mem[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12341_ (.D(_00220_),
    .CLK(clknet_leaf_79_clock),
    .Q(\u2.mem[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12342_ (.D(_00221_),
    .CLK(clknet_leaf_78_clock),
    .Q(\u2.mem[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12343_ (.D(_00222_),
    .CLK(clknet_leaf_132_clock),
    .Q(\u2.mem[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12344_ (.D(_00223_),
    .CLK(clknet_leaf_131_clock),
    .Q(\u2.mem[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12345_ (.D(_00224_),
    .CLK(clknet_leaf_60_clock),
    .Q(\u2.mem[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12346_ (.D(_00225_),
    .CLK(clknet_leaf_59_clock),
    .Q(\u2.mem[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12347_ (.D(_00226_),
    .CLK(clknet_leaf_221_clock),
    .Q(\u2.mem[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12348_ (.D(_00227_),
    .CLK(clknet_leaf_202_clock),
    .Q(\u2.mem[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12349_ (.D(_00228_),
    .CLK(clknet_leaf_202_clock),
    .Q(\u2.mem[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12350_ (.D(_00229_),
    .CLK(clknet_leaf_201_clock),
    .Q(\u2.mem[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12351_ (.D(_00230_),
    .CLK(clknet_leaf_148_clock),
    .Q(\u2.mem[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12352_ (.D(_00231_),
    .CLK(clknet_leaf_148_clock),
    .Q(\u2.mem[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12353_ (.D(_00232_),
    .CLK(clknet_leaf_150_clock),
    .Q(\u2.mem[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12354_ (.D(_00233_),
    .CLK(clknet_leaf_150_clock),
    .Q(\u2.mem[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12355_ (.D(_00234_),
    .CLK(clknet_leaf_83_clock),
    .Q(\u2.mem[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12356_ (.D(_00235_),
    .CLK(clknet_leaf_80_clock),
    .Q(\u2.mem[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12357_ (.D(_00236_),
    .CLK(clknet_leaf_80_clock),
    .Q(\u2.mem[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12358_ (.D(_00237_),
    .CLK(clknet_leaf_80_clock),
    .Q(\u2.mem[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12359_ (.D(_00238_),
    .CLK(clknet_leaf_133_clock),
    .Q(\u2.mem[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12360_ (.D(_00239_),
    .CLK(clknet_leaf_136_clock),
    .Q(\u2.mem[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12361_ (.D(_00240_),
    .CLK(clknet_leaf_133_clock),
    .Q(\u2.mem[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12362_ (.D(_00241_),
    .CLK(clknet_leaf_134_clock),
    .Q(\u2.mem[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12363_ (.D(_00242_),
    .CLK(clknet_leaf_208_clock),
    .Q(\u2.mem[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12364_ (.D(_00243_),
    .CLK(clknet_leaf_206_clock),
    .Q(\u2.mem[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12365_ (.D(_00244_),
    .CLK(clknet_leaf_210_clock),
    .Q(\u2.mem[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12366_ (.D(_00245_),
    .CLK(clknet_leaf_209_clock),
    .Q(\u2.mem[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12367_ (.D(_00246_),
    .CLK(clknet_leaf_223_clock),
    .Q(\u2.mem[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12368_ (.D(_00247_),
    .CLK(clknet_leaf_222_clock),
    .Q(\u2.mem[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12369_ (.D(_00248_),
    .CLK(clknet_leaf_223_clock),
    .Q(\u2.mem[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12370_ (.D(_00249_),
    .CLK(clknet_leaf_150_clock),
    .Q(\u2.mem[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12371_ (.D(_00250_),
    .CLK(clknet_leaf_78_clock),
    .Q(\u2.mem[15][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12372_ (.D(_00251_),
    .CLK(clknet_leaf_80_clock),
    .Q(\u2.mem[15][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12373_ (.D(_00252_),
    .CLK(clknet_leaf_79_clock),
    .Q(\u2.mem[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12374_ (.D(_00253_),
    .CLK(clknet_leaf_78_clock),
    .Q(\u2.mem[15][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12375_ (.D(_00254_),
    .CLK(clknet_leaf_59_clock),
    .Q(\u2.mem[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12376_ (.D(_00255_),
    .CLK(clknet_leaf_131_clock),
    .Q(\u2.mem[15][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12377_ (.D(_00256_),
    .CLK(clknet_leaf_60_clock),
    .Q(\u2.mem[15][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12378_ (.D(_00257_),
    .CLK(clknet_leaf_60_clock),
    .Q(\u2.mem[15][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12379_ (.D(_00258_),
    .CLK(clknet_leaf_207_clock),
    .Q(\u2.mem[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12380_ (.D(_00259_),
    .CLK(clknet_leaf_205_clock),
    .Q(\u2.mem[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12381_ (.D(_00260_),
    .CLK(clknet_leaf_206_clock),
    .Q(\u2.mem[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12382_ (.D(_00261_),
    .CLK(clknet_leaf_207_clock),
    .Q(\u2.mem[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12383_ (.D(_00262_),
    .CLK(clknet_leaf_223_clock),
    .Q(\u2.mem[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12384_ (.D(_00263_),
    .CLK(clknet_leaf_221_clock),
    .Q(\u2.mem[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12385_ (.D(_00264_),
    .CLK(clknet_leaf_223_clock),
    .Q(\u2.mem[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12386_ (.D(_00265_),
    .CLK(clknet_leaf_224_clock),
    .Q(\u2.mem[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12387_ (.D(_00266_),
    .CLK(clknet_leaf_77_clock),
    .Q(\u2.mem[16][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12388_ (.D(_00267_),
    .CLK(clknet_leaf_81_clock),
    .Q(\u2.mem[16][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12389_ (.D(_00268_),
    .CLK(clknet_leaf_78_clock),
    .Q(\u2.mem[16][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12390_ (.D(_00269_),
    .CLK(clknet_leaf_77_clock),
    .Q(\u2.mem[16][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12391_ (.D(_00270_),
    .CLK(clknet_leaf_134_clock),
    .Q(\u2.mem[16][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12392_ (.D(_00271_),
    .CLK(clknet_leaf_133_clock),
    .Q(\u2.mem[16][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12393_ (.D(_00272_),
    .CLK(clknet_leaf_132_clock),
    .Q(\u2.mem[16][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12394_ (.D(_00273_),
    .CLK(clknet_leaf_134_clock),
    .Q(\u2.mem[16][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12395_ (.D(_00274_),
    .CLK(clknet_leaf_179_clock),
    .Q(\u2.mem[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12396_ (.D(_00275_),
    .CLK(clknet_leaf_180_clock),
    .Q(\u2.mem[17][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12397_ (.D(_00276_),
    .CLK(clknet_leaf_180_clock),
    .Q(\u2.mem[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12398_ (.D(_00277_),
    .CLK(clknet_leaf_179_clock),
    .Q(\u2.mem[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12399_ (.D(_00278_),
    .CLK(clknet_leaf_155_clock),
    .Q(\u2.mem[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12400_ (.D(_00279_),
    .CLK(clknet_leaf_156_clock),
    .Q(\u2.mem[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12401_ (.D(_00280_),
    .CLK(clknet_leaf_161_clock),
    .Q(\u2.mem[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12402_ (.D(_00281_),
    .CLK(clknet_leaf_155_clock),
    .Q(\u2.mem[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12403_ (.D(_00282_),
    .CLK(clknet_leaf_108_clock),
    .Q(\u2.mem[17][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12404_ (.D(_00283_),
    .CLK(clknet_leaf_107_clock),
    .Q(\u2.mem[17][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12405_ (.D(_00284_),
    .CLK(clknet_leaf_88_clock),
    .Q(\u2.mem[17][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12406_ (.D(_00285_),
    .CLK(clknet_leaf_88_clock),
    .Q(\u2.mem[17][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12407_ (.D(_00286_),
    .CLK(clknet_leaf_112_clock),
    .Q(\u2.mem[17][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12408_ (.D(_00287_),
    .CLK(clknet_leaf_122_clock),
    .Q(\u2.mem[17][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12409_ (.D(_00288_),
    .CLK(clknet_leaf_122_clock),
    .Q(\u2.mem[17][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12410_ (.D(_00289_),
    .CLK(clknet_leaf_112_clock),
    .Q(\u2.mem[17][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12411_ (.D(_00290_),
    .CLK(clknet_leaf_177_clock),
    .Q(\u2.mem[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12412_ (.D(_00291_),
    .CLK(clknet_leaf_198_clock),
    .Q(\u2.mem[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12413_ (.D(_00292_),
    .CLK(clknet_leaf_197_clock),
    .Q(\u2.mem[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12414_ (.D(_00293_),
    .CLK(clknet_leaf_178_clock),
    .Q(\u2.mem[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12415_ (.D(_00294_),
    .CLK(clknet_leaf_160_clock),
    .Q(\u2.mem[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12416_ (.D(_00295_),
    .CLK(clknet_leaf_160_clock),
    .Q(\u2.mem[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12417_ (.D(_00296_),
    .CLK(clknet_leaf_161_clock),
    .Q(\u2.mem[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12418_ (.D(_00297_),
    .CLK(clknet_leaf_160_clock),
    .Q(\u2.mem[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12419_ (.D(_00298_),
    .CLK(clknet_leaf_110_clock),
    .Q(\u2.mem[18][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12420_ (.D(_00299_),
    .CLK(clknet_leaf_108_clock),
    .Q(\u2.mem[18][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12421_ (.D(_00300_),
    .CLK(clknet_leaf_87_clock),
    .Q(\u2.mem[18][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12422_ (.D(_00301_),
    .CLK(clknet_leaf_87_clock),
    .Q(\u2.mem[18][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12423_ (.D(_00302_),
    .CLK(clknet_leaf_128_clock),
    .Q(\u2.mem[18][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12424_ (.D(_00303_),
    .CLK(clknet_leaf_123_clock),
    .Q(\u2.mem[18][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12425_ (.D(_00304_),
    .CLK(clknet_leaf_128_clock),
    .Q(\u2.mem[18][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12426_ (.D(_00305_),
    .CLK(clknet_leaf_112_clock),
    .Q(\u2.mem[18][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12427_ (.D(_00306_),
    .CLK(clknet_leaf_178_clock),
    .Q(\u2.mem[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12428_ (.D(_00307_),
    .CLK(clknet_leaf_180_clock),
    .Q(\u2.mem[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12429_ (.D(_00308_),
    .CLK(clknet_leaf_196_clock),
    .Q(\u2.mem[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12430_ (.D(_00309_),
    .CLK(clknet_leaf_178_clock),
    .Q(\u2.mem[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12431_ (.D(_00310_),
    .CLK(clknet_leaf_160_clock),
    .Q(\u2.mem[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12432_ (.D(_00311_),
    .CLK(clknet_leaf_159_clock),
    .Q(\u2.mem[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12433_ (.D(_00312_),
    .CLK(clknet_leaf_161_clock),
    .Q(\u2.mem[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12434_ (.D(_00313_),
    .CLK(clknet_leaf_124_clock),
    .Q(\u2.mem[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12435_ (.D(_00314_),
    .CLK(clknet_leaf_108_clock),
    .Q(\u2.mem[19][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12436_ (.D(_00315_),
    .CLK(clknet_leaf_107_clock),
    .Q(\u2.mem[19][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12437_ (.D(_00316_),
    .CLK(clknet_leaf_88_clock),
    .Q(\u2.mem[19][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12438_ (.D(_00317_),
    .CLK(clknet_leaf_87_clock),
    .Q(\u2.mem[19][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12439_ (.D(_00318_),
    .CLK(clknet_leaf_127_clock),
    .Q(\u2.mem[19][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12440_ (.D(_00319_),
    .CLK(clknet_leaf_123_clock),
    .Q(\u2.mem[19][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12441_ (.D(_00320_),
    .CLK(clknet_leaf_127_clock),
    .Q(\u2.mem[19][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12442_ (.D(_00321_),
    .CLK(clknet_leaf_128_clock),
    .Q(\u2.mem[19][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12443_ (.D(_00322_),
    .CLK(clknet_leaf_199_clock),
    .Q(\u2.mem[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12444_ (.D(_00323_),
    .CLK(clknet_leaf_198_clock),
    .Q(\u2.mem[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12445_ (.D(_00324_),
    .CLK(clknet_leaf_198_clock),
    .Q(\u2.mem[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12446_ (.D(_00325_),
    .CLK(clknet_leaf_199_clock),
    .Q(\u2.mem[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12447_ (.D(_00326_),
    .CLK(clknet_leaf_159_clock),
    .Q(\u2.mem[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12448_ (.D(_00327_),
    .CLK(clknet_leaf_159_clock),
    .Q(\u2.mem[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12449_ (.D(_00328_),
    .CLK(clknet_leaf_159_clock),
    .Q(\u2.mem[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12450_ (.D(_00329_),
    .CLK(clknet_leaf_159_clock),
    .Q(\u2.mem[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12451_ (.D(_00330_),
    .CLK(clknet_leaf_84_clock),
    .Q(\u2.mem[20][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12452_ (.D(_00331_),
    .CLK(clknet_leaf_84_clock),
    .Q(\u2.mem[20][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12453_ (.D(_00332_),
    .CLK(clknet_leaf_86_clock),
    .Q(\u2.mem[20][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12454_ (.D(_00333_),
    .CLK(clknet_leaf_85_clock),
    .Q(\u2.mem[20][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12455_ (.D(_00334_),
    .CLK(clknet_leaf_127_clock),
    .Q(\u2.mem[20][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12456_ (.D(_00335_),
    .CLK(clknet_leaf_126_clock),
    .Q(\u2.mem[20][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12457_ (.D(_00336_),
    .CLK(clknet_leaf_126_clock),
    .Q(\u2.mem[20][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12458_ (.D(_00337_),
    .CLK(clknet_leaf_127_clock),
    .Q(\u2.mem[20][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12459_ (.D(_00338_),
    .CLK(clknet_leaf_179_clock),
    .Q(\u2.mem[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12460_ (.D(_00339_),
    .CLK(clknet_leaf_196_clock),
    .Q(\u2.mem[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12461_ (.D(_00340_),
    .CLK(clknet_leaf_196_clock),
    .Q(\u2.mem[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12462_ (.D(_00341_),
    .CLK(clknet_leaf_191_clock),
    .Q(\u2.mem[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12463_ (.D(_00342_),
    .CLK(clknet_leaf_172_clock),
    .Q(\u2.mem[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12464_ (.D(_00343_),
    .CLK(clknet_leaf_173_clock),
    .Q(\u2.mem[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12465_ (.D(_00344_),
    .CLK(clknet_leaf_167_clock),
    .Q(\u2.mem[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12466_ (.D(_00345_),
    .CLK(clknet_leaf_162_clock),
    .Q(\u2.mem[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12467_ (.D(_00346_),
    .CLK(clknet_leaf_108_clock),
    .Q(\u2.mem[21][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12468_ (.D(_00347_),
    .CLK(clknet_leaf_105_clock),
    .Q(\u2.mem[21][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12469_ (.D(_00348_),
    .CLK(clknet_leaf_106_clock),
    .Q(\u2.mem[21][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12470_ (.D(_00349_),
    .CLK(clknet_leaf_106_clock),
    .Q(\u2.mem[21][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12471_ (.D(_00350_),
    .CLK(clknet_leaf_122_clock),
    .Q(\u2.mem[21][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12472_ (.D(_00351_),
    .CLK(clknet_leaf_121_clock),
    .Q(\u2.mem[21][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12473_ (.D(_00352_),
    .CLK(clknet_leaf_122_clock),
    .Q(\u2.mem[21][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12474_ (.D(_00353_),
    .CLK(clknet_leaf_123_clock),
    .Q(\u2.mem[21][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12475_ (.D(_00354_),
    .CLK(clknet_leaf_182_clock),
    .Q(\u2.mem[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12476_ (.D(_00355_),
    .CLK(clknet_leaf_181_clock),
    .Q(\u2.mem[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12477_ (.D(_00356_),
    .CLK(clknet_leaf_181_clock),
    .Q(\u2.mem[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12478_ (.D(_00357_),
    .CLK(clknet_leaf_181_clock),
    .Q(\u2.mem[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12479_ (.D(_00358_),
    .CLK(clknet_leaf_163_clock),
    .Q(\u2.mem[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12480_ (.D(_00359_),
    .CLK(clknet_leaf_164_clock),
    .Q(\u2.mem[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12481_ (.D(_00360_),
    .CLK(clknet_leaf_164_clock),
    .Q(\u2.mem[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12482_ (.D(_00361_),
    .CLK(clknet_leaf_164_clock),
    .Q(\u2.mem[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12483_ (.D(_00362_),
    .CLK(clknet_leaf_123_clock),
    .Q(\u2.mem[22][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12484_ (.D(_00363_),
    .CLK(clknet_leaf_105_clock),
    .Q(\u2.mem[22][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12485_ (.D(_00364_),
    .CLK(clknet_leaf_100_clock),
    .Q(\u2.mem[22][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12486_ (.D(_00365_),
    .CLK(clknet_leaf_100_clock),
    .Q(\u2.mem[22][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12487_ (.D(_00366_),
    .CLK(clknet_leaf_121_clock),
    .Q(\u2.mem[22][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12488_ (.D(_00367_),
    .CLK(clknet_leaf_164_clock),
    .Q(\u2.mem[22][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12489_ (.D(_00368_),
    .CLK(clknet_leaf_121_clock),
    .Q(\u2.mem[22][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12490_ (.D(_00369_),
    .CLK(clknet_leaf_121_clock),
    .Q(\u2.mem[22][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12491_ (.D(_00370_),
    .CLK(clknet_leaf_182_clock),
    .Q(\u2.mem[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12492_ (.D(_00371_),
    .CLK(clknet_leaf_190_clock),
    .Q(\u2.mem[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12493_ (.D(_00372_),
    .CLK(clknet_leaf_186_clock),
    .Q(\u2.mem[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12494_ (.D(_00373_),
    .CLK(clknet_leaf_181_clock),
    .Q(\u2.mem[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12495_ (.D(_00374_),
    .CLK(clknet_leaf_163_clock),
    .Q(\u2.mem[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12496_ (.D(_00375_),
    .CLK(clknet_leaf_163_clock),
    .Q(\u2.mem[23][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12497_ (.D(_00376_),
    .CLK(clknet_leaf_163_clock),
    .Q(\u2.mem[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12498_ (.D(_00377_),
    .CLK(clknet_leaf_161_clock),
    .Q(\u2.mem[23][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12499_ (.D(_00378_),
    .CLK(clknet_leaf_123_clock),
    .Q(\u2.mem[23][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12500_ (.D(_00379_),
    .CLK(clknet_leaf_105_clock),
    .Q(\u2.mem[23][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12501_ (.D(_00380_),
    .CLK(clknet_leaf_106_clock),
    .Q(\u2.mem[23][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12502_ (.D(_00381_),
    .CLK(clknet_leaf_106_clock),
    .Q(\u2.mem[23][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12503_ (.D(_00382_),
    .CLK(clknet_leaf_121_clock),
    .Q(\u2.mem[23][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12504_ (.D(_00383_),
    .CLK(clknet_leaf_121_clock),
    .Q(\u2.mem[23][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12505_ (.D(_00384_),
    .CLK(clknet_leaf_163_clock),
    .Q(\u2.mem[23][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12506_ (.D(_00385_),
    .CLK(clknet_leaf_121_clock),
    .Q(\u2.mem[23][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12507_ (.D(_00386_),
    .CLK(clknet_leaf_179_clock),
    .Q(\u2.mem[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12508_ (.D(_00387_),
    .CLK(clknet_leaf_180_clock),
    .Q(\u2.mem[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12509_ (.D(_00388_),
    .CLK(clknet_leaf_180_clock),
    .Q(\u2.mem[24][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12510_ (.D(_00389_),
    .CLK(clknet_leaf_179_clock),
    .Q(\u2.mem[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12511_ (.D(_00390_),
    .CLK(clknet_leaf_162_clock),
    .Q(\u2.mem[24][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12512_ (.D(_00391_),
    .CLK(clknet_leaf_162_clock),
    .Q(\u2.mem[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12513_ (.D(_00392_),
    .CLK(clknet_leaf_162_clock),
    .Q(\u2.mem[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12514_ (.D(_00393_),
    .CLK(clknet_leaf_162_clock),
    .Q(\u2.mem[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12515_ (.D(_00394_),
    .CLK(clknet_leaf_105_clock),
    .Q(\u2.mem[24][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12516_ (.D(_00395_),
    .CLK(clknet_leaf_99_clock),
    .Q(\u2.mem[24][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12517_ (.D(_00396_),
    .CLK(clknet_leaf_95_clock),
    .Q(\u2.mem[24][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12518_ (.D(_00397_),
    .CLK(clknet_leaf_94_clock),
    .Q(\u2.mem[24][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12519_ (.D(_00398_),
    .CLK(clknet_leaf_117_clock),
    .Q(\u2.mem[24][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12520_ (.D(_00399_),
    .CLK(clknet_leaf_118_clock),
    .Q(\u2.mem[24][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12521_ (.D(_00400_),
    .CLK(clknet_leaf_118_clock),
    .Q(\u2.mem[24][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12522_ (.D(_00401_),
    .CLK(clknet_leaf_112_clock),
    .Q(\u2.mem[24][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12523_ (.D(_00402_),
    .CLK(clknet_leaf_183_clock),
    .Q(\u2.mem[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12524_ (.D(_00403_),
    .CLK(clknet_leaf_187_clock),
    .Q(\u2.mem[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12525_ (.D(_00404_),
    .CLK(clknet_leaf_188_clock),
    .Q(\u2.mem[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12526_ (.D(_00405_),
    .CLK(clknet_leaf_187_clock),
    .Q(\u2.mem[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12527_ (.D(_00406_),
    .CLK(clknet_leaf_169_clock),
    .Q(\u2.mem[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12528_ (.D(_00407_),
    .CLK(clknet_leaf_169_clock),
    .Q(\u2.mem[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12529_ (.D(_00408_),
    .CLK(clknet_leaf_166_clock),
    .Q(\u2.mem[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12530_ (.D(_00409_),
    .CLK(clknet_leaf_166_clock),
    .Q(\u2.mem[25][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12531_ (.D(_00410_),
    .CLK(clknet_leaf_103_clock),
    .Q(\u2.mem[25][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12532_ (.D(_00411_),
    .CLK(clknet_leaf_98_clock),
    .Q(\u2.mem[25][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12533_ (.D(_00412_),
    .CLK(clknet_leaf_98_clock),
    .Q(\u2.mem[25][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12534_ (.D(_00413_),
    .CLK(clknet_leaf_97_clock),
    .Q(\u2.mem[25][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12535_ (.D(_00414_),
    .CLK(clknet_leaf_115_clock),
    .Q(\u2.mem[25][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12536_ (.D(_00415_),
    .CLK(clknet_leaf_116_clock),
    .Q(\u2.mem[25][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12537_ (.D(_00416_),
    .CLK(clknet_leaf_116_clock),
    .Q(\u2.mem[25][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12538_ (.D(_00417_),
    .CLK(clknet_leaf_115_clock),
    .Q(\u2.mem[25][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12539_ (.D(_00418_),
    .CLK(clknet_leaf_184_clock),
    .Q(\u2.mem[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12540_ (.D(_00419_),
    .CLK(clknet_leaf_189_clock),
    .Q(\u2.mem[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12541_ (.D(_00420_),
    .CLK(clknet_leaf_188_clock),
    .Q(\u2.mem[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12542_ (.D(_00421_),
    .CLK(clknet_leaf_188_clock),
    .Q(\u2.mem[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12543_ (.D(_00422_),
    .CLK(clknet_leaf_168_clock),
    .Q(\u2.mem[26][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12544_ (.D(_00423_),
    .CLK(clknet_leaf_168_clock),
    .Q(\u2.mem[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12545_ (.D(_00424_),
    .CLK(clknet_leaf_168_clock),
    .Q(\u2.mem[26][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12546_ (.D(_00425_),
    .CLK(clknet_leaf_168_clock),
    .Q(\u2.mem[26][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12547_ (.D(_00426_),
    .CLK(clknet_leaf_103_clock),
    .Q(\u2.mem[26][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12548_ (.D(_00427_),
    .CLK(clknet_leaf_98_clock),
    .Q(\u2.mem[26][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12549_ (.D(_00428_),
    .CLK(clknet_leaf_98_clock),
    .Q(\u2.mem[26][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12550_ (.D(_00429_),
    .CLK(clknet_leaf_98_clock),
    .Q(\u2.mem[26][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12551_ (.D(_00430_),
    .CLK(clknet_leaf_115_clock),
    .Q(\u2.mem[26][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12552_ (.D(_00431_),
    .CLK(clknet_leaf_119_clock),
    .Q(\u2.mem[26][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12553_ (.D(_00432_),
    .CLK(clknet_leaf_119_clock),
    .Q(\u2.mem[26][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12554_ (.D(_00433_),
    .CLK(clknet_leaf_119_clock),
    .Q(\u2.mem[26][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12555_ (.D(_00434_),
    .CLK(clknet_leaf_191_clock),
    .Q(\u2.mem[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12556_ (.D(_00435_),
    .CLK(clknet_leaf_190_clock),
    .Q(\u2.mem[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12557_ (.D(_00436_),
    .CLK(clknet_leaf_192_clock),
    .Q(\u2.mem[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12558_ (.D(_00437_),
    .CLK(clknet_leaf_191_clock),
    .Q(\u2.mem[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12559_ (.D(_00438_),
    .CLK(clknet_leaf_170_clock),
    .Q(\u2.mem[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12560_ (.D(_00439_),
    .CLK(clknet_leaf_171_clock),
    .Q(\u2.mem[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12561_ (.D(_00440_),
    .CLK(clknet_leaf_170_clock),
    .Q(\u2.mem[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12562_ (.D(_00441_),
    .CLK(clknet_leaf_171_clock),
    .Q(\u2.mem[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12563_ (.D(_00442_),
    .CLK(clknet_leaf_94_clock),
    .Q(\u2.mem[27][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12564_ (.D(_00443_),
    .CLK(clknet_leaf_95_clock),
    .Q(\u2.mem[27][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12565_ (.D(_00444_),
    .CLK(clknet_leaf_96_clock),
    .Q(\u2.mem[27][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12566_ (.D(_00445_),
    .CLK(clknet_leaf_94_clock),
    .Q(\u2.mem[27][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12567_ (.D(_00446_),
    .CLK(clknet_leaf_113_clock),
    .Q(\u2.mem[27][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12568_ (.D(_00447_),
    .CLK(clknet_leaf_112_clock),
    .Q(\u2.mem[27][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12569_ (.D(_00448_),
    .CLK(clknet_leaf_113_clock),
    .Q(\u2.mem[27][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12570_ (.D(_00449_),
    .CLK(clknet_leaf_111_clock),
    .Q(\u2.mem[27][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12571_ (.D(_00450_),
    .CLK(clknet_leaf_182_clock),
    .Q(\u2.mem[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12572_ (.D(_00451_),
    .CLK(clknet_leaf_186_clock),
    .Q(\u2.mem[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12573_ (.D(_00452_),
    .CLK(clknet_leaf_187_clock),
    .Q(\u2.mem[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12574_ (.D(_00453_),
    .CLK(clknet_leaf_186_clock),
    .Q(\u2.mem[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12575_ (.D(_00454_),
    .CLK(clknet_leaf_183_clock),
    .Q(\u2.mem[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12576_ (.D(_00455_),
    .CLK(clknet_leaf_169_clock),
    .Q(\u2.mem[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12577_ (.D(_00456_),
    .CLK(clknet_leaf_170_clock),
    .Q(\u2.mem[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12578_ (.D(_00457_),
    .CLK(clknet_leaf_169_clock),
    .Q(\u2.mem[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12579_ (.D(_00458_),
    .CLK(clknet_leaf_104_clock),
    .Q(\u2.mem[28][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12580_ (.D(_00459_),
    .CLK(clknet_leaf_98_clock),
    .Q(\u2.mem[28][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12581_ (.D(_00460_),
    .CLK(clknet_leaf_98_clock),
    .Q(\u2.mem[28][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12582_ (.D(_00461_),
    .CLK(clknet_leaf_100_clock),
    .Q(\u2.mem[28][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12583_ (.D(_00462_),
    .CLK(clknet_leaf_115_clock),
    .Q(\u2.mem[28][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12584_ (.D(_00463_),
    .CLK(clknet_leaf_115_clock),
    .Q(\u2.mem[28][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12585_ (.D(_00464_),
    .CLK(clknet_leaf_115_clock),
    .Q(\u2.mem[28][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12586_ (.D(_00465_),
    .CLK(clknet_leaf_115_clock),
    .Q(\u2.mem[28][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12587_ (.D(_00466_),
    .CLK(clknet_leaf_186_clock),
    .Q(\u2.mem[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12588_ (.D(_00467_),
    .CLK(clknet_leaf_190_clock),
    .Q(\u2.mem[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12589_ (.D(_00468_),
    .CLK(clknet_leaf_187_clock),
    .Q(\u2.mem[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12590_ (.D(_00469_),
    .CLK(clknet_leaf_190_clock),
    .Q(\u2.mem[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12591_ (.D(_00470_),
    .CLK(clknet_leaf_172_clock),
    .Q(\u2.mem[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12592_ (.D(_00471_),
    .CLK(clknet_leaf_168_clock),
    .Q(\u2.mem[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12593_ (.D(_00472_),
    .CLK(clknet_leaf_167_clock),
    .Q(\u2.mem[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12594_ (.D(_00473_),
    .CLK(clknet_leaf_167_clock),
    .Q(\u2.mem[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12595_ (.D(_00474_),
    .CLK(clknet_leaf_105_clock),
    .Q(\u2.mem[29][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12596_ (.D(_00475_),
    .CLK(clknet_leaf_99_clock),
    .Q(\u2.mem[29][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12597_ (.D(_00476_),
    .CLK(clknet_leaf_99_clock),
    .Q(\u2.mem[29][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12598_ (.D(_00477_),
    .CLK(clknet_leaf_96_clock),
    .Q(\u2.mem[29][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12599_ (.D(_00478_),
    .CLK(clknet_leaf_113_clock),
    .Q(\u2.mem[29][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12600_ (.D(_00479_),
    .CLK(clknet_leaf_117_clock),
    .Q(\u2.mem[29][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12601_ (.D(_00480_),
    .CLK(clknet_leaf_116_clock),
    .Q(\u2.mem[29][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12602_ (.D(_00481_),
    .CLK(clknet_leaf_113_clock),
    .Q(\u2.mem[29][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12603_ (.D(_00482_),
    .CLK(clknet_leaf_196_clock),
    .Q(\u2.mem[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12604_ (.D(_00483_),
    .CLK(clknet_leaf_191_clock),
    .Q(\u2.mem[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12605_ (.D(_00484_),
    .CLK(clknet_leaf_196_clock),
    .Q(\u2.mem[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12606_ (.D(_00485_),
    .CLK(clknet_leaf_195_clock),
    .Q(\u2.mem[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12607_ (.D(_00486_),
    .CLK(clknet_leaf_173_clock),
    .Q(\u2.mem[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12608_ (.D(_00487_),
    .CLK(clknet_leaf_172_clock),
    .Q(\u2.mem[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12609_ (.D(_00488_),
    .CLK(clknet_leaf_155_clock),
    .Q(\u2.mem[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12610_ (.D(_00489_),
    .CLK(clknet_leaf_173_clock),
    .Q(\u2.mem[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12611_ (.D(_00490_),
    .CLK(clknet_leaf_94_clock),
    .Q(\u2.mem[30][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12612_ (.D(_00491_),
    .CLK(clknet_leaf_93_clock),
    .Q(\u2.mem[30][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12613_ (.D(_00492_),
    .CLK(clknet_leaf_94_clock),
    .Q(\u2.mem[30][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12614_ (.D(_00493_),
    .CLK(clknet_leaf_93_clock),
    .Q(\u2.mem[30][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12615_ (.D(_00494_),
    .CLK(clknet_leaf_113_clock),
    .Q(\u2.mem[30][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12616_ (.D(_00495_),
    .CLK(clknet_leaf_113_clock),
    .Q(\u2.mem[30][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12617_ (.D(_00496_),
    .CLK(clknet_leaf_111_clock),
    .Q(\u2.mem[30][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12618_ (.D(_00497_),
    .CLK(clknet_leaf_111_clock),
    .Q(\u2.mem[30][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12619_ (.D(_00498_),
    .CLK(clknet_leaf_186_clock),
    .Q(\u2.mem[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12620_ (.D(_00499_),
    .CLK(clknet_leaf_190_clock),
    .Q(\u2.mem[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12621_ (.D(_00500_),
    .CLK(clknet_leaf_190_clock),
    .Q(\u2.mem[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12622_ (.D(_00501_),
    .CLK(clknet_leaf_189_clock),
    .Q(\u2.mem[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12623_ (.D(_00502_),
    .CLK(clknet_leaf_172_clock),
    .Q(\u2.mem[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12624_ (.D(_00503_),
    .CLK(clknet_leaf_168_clock),
    .Q(\u2.mem[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12625_ (.D(_00504_),
    .CLK(clknet_leaf_172_clock),
    .Q(\u2.mem[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12626_ (.D(_00505_),
    .CLK(clknet_leaf_170_clock),
    .Q(\u2.mem[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12627_ (.D(_00506_),
    .CLK(clknet_leaf_97_clock),
    .Q(\u2.mem[31][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12628_ (.D(_00507_),
    .CLK(clknet_leaf_97_clock),
    .Q(\u2.mem[31][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12629_ (.D(_00508_),
    .CLK(clknet_leaf_97_clock),
    .Q(\u2.mem[31][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12630_ (.D(_00509_),
    .CLK(clknet_leaf_96_clock),
    .Q(\u2.mem[31][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12631_ (.D(_00510_),
    .CLK(clknet_leaf_114_clock),
    .Q(\u2.mem[31][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12632_ (.D(_00511_),
    .CLK(clknet_leaf_104_clock),
    .Q(\u2.mem[31][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12633_ (.D(_00512_),
    .CLK(clknet_leaf_103_clock),
    .Q(\u2.mem[31][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12634_ (.D(_00513_),
    .CLK(clknet_leaf_114_clock),
    .Q(\u2.mem[31][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12635_ (.D(_00514_),
    .CLK(clknet_leaf_194_clock),
    .Q(\u2.mem[32][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12636_ (.D(_00515_),
    .CLK(clknet_leaf_192_clock),
    .Q(\u2.mem[32][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12637_ (.D(_00516_),
    .CLK(clknet_leaf_192_clock),
    .Q(\u2.mem[32][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12638_ (.D(_00517_),
    .CLK(clknet_leaf_192_clock),
    .Q(\u2.mem[32][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12639_ (.D(_00518_),
    .CLK(clknet_leaf_175_clock),
    .Q(\u2.mem[32][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12640_ (.D(_00519_),
    .CLK(clknet_leaf_172_clock),
    .Q(\u2.mem[32][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12641_ (.D(_00520_),
    .CLK(clknet_leaf_173_clock),
    .Q(\u2.mem[32][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12642_ (.D(_00521_),
    .CLK(clknet_leaf_174_clock),
    .Q(\u2.mem[32][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12643_ (.D(_00522_),
    .CLK(clknet_leaf_94_clock),
    .Q(\u2.mem[32][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12644_ (.D(_00523_),
    .CLK(clknet_leaf_92_clock),
    .Q(\u2.mem[32][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12645_ (.D(_00524_),
    .CLK(clknet_leaf_93_clock),
    .Q(\u2.mem[32][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12646_ (.D(_00525_),
    .CLK(clknet_leaf_93_clock),
    .Q(\u2.mem[32][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12647_ (.D(_00526_),
    .CLK(clknet_leaf_114_clock),
    .Q(\u2.mem[32][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12648_ (.D(_00527_),
    .CLK(clknet_leaf_114_clock),
    .Q(\u2.mem[32][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12649_ (.D(_00528_),
    .CLK(clknet_leaf_111_clock),
    .Q(\u2.mem[32][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12650_ (.D(_00529_),
    .CLK(clknet_leaf_110_clock),
    .Q(\u2.mem[32][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12651_ (.D(_00530_),
    .CLK(clknet_leaf_207_clock),
    .Q(\u2.mem[33][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12652_ (.D(_00531_),
    .CLK(clknet_leaf_205_clock),
    .Q(\u2.mem[33][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12653_ (.D(_00532_),
    .CLK(clknet_leaf_205_clock),
    .Q(\u2.mem[33][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12654_ (.D(_00533_),
    .CLK(clknet_leaf_205_clock),
    .Q(\u2.mem[33][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12655_ (.D(_00534_),
    .CLK(clknet_leaf_223_clock),
    .Q(\u2.mem[33][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12656_ (.D(_00535_),
    .CLK(clknet_leaf_221_clock),
    .Q(\u2.mem[33][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12657_ (.D(_00536_),
    .CLK(clknet_leaf_224_clock),
    .Q(\u2.mem[33][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12658_ (.D(_00537_),
    .CLK(clknet_leaf_224_clock),
    .Q(\u2.mem[33][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12659_ (.D(_00538_),
    .CLK(clknet_leaf_81_clock),
    .Q(\u2.mem[33][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12660_ (.D(_00539_),
    .CLK(clknet_leaf_75_clock),
    .Q(\u2.mem[33][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12661_ (.D(_00540_),
    .CLK(clknet_leaf_77_clock),
    .Q(\u2.mem[33][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12662_ (.D(_00541_),
    .CLK(clknet_leaf_76_clock),
    .Q(\u2.mem[33][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12663_ (.D(_00542_),
    .CLK(clknet_leaf_58_clock),
    .Q(\u2.mem[33][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12664_ (.D(_00543_),
    .CLK(clknet_leaf_135_clock),
    .Q(\u2.mem[33][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12665_ (.D(_00544_),
    .CLK(clknet_leaf_58_clock),
    .Q(\u2.mem[33][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12666_ (.D(_00545_),
    .CLK(clknet_leaf_56_clock),
    .Q(\u2.mem[33][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12667_ (.D(_00546_),
    .CLK(clknet_leaf_195_clock),
    .Q(\u2.mem[34][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12668_ (.D(_00547_),
    .CLK(clknet_leaf_193_clock),
    .Q(\u2.mem[34][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12669_ (.D(_00548_),
    .CLK(clknet_leaf_193_clock),
    .Q(\u2.mem[34][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12670_ (.D(_00549_),
    .CLK(clknet_leaf_194_clock),
    .Q(\u2.mem[34][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12671_ (.D(_00550_),
    .CLK(clknet_leaf_177_clock),
    .Q(\u2.mem[34][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12672_ (.D(_00551_),
    .CLK(clknet_leaf_177_clock),
    .Q(\u2.mem[34][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12673_ (.D(_00552_),
    .CLK(clknet_leaf_154_clock),
    .Q(\u2.mem[34][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12674_ (.D(_00553_),
    .CLK(clknet_leaf_154_clock),
    .Q(\u2.mem[34][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12675_ (.D(_00554_),
    .CLK(clknet_leaf_86_clock),
    .Q(\u2.mem[34][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12676_ (.D(_00555_),
    .CLK(clknet_leaf_90_clock),
    .Q(\u2.mem[34][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12677_ (.D(_00556_),
    .CLK(clknet_leaf_90_clock),
    .Q(\u2.mem[34][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12678_ (.D(_00557_),
    .CLK(clknet_leaf_89_clock),
    .Q(\u2.mem[34][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12679_ (.D(_00558_),
    .CLK(clknet_leaf_130_clock),
    .Q(\u2.mem[34][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12680_ (.D(_00559_),
    .CLK(clknet_leaf_129_clock),
    .Q(\u2.mem[34][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12681_ (.D(_00560_),
    .CLK(clknet_leaf_129_clock),
    .Q(\u2.mem[34][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12682_ (.D(_00561_),
    .CLK(clknet_leaf_127_clock),
    .Q(\u2.mem[34][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12683_ (.D(_00562_),
    .CLK(clknet_leaf_195_clock),
    .Q(\u2.mem[35][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12684_ (.D(_00563_),
    .CLK(clknet_leaf_193_clock),
    .Q(\u2.mem[35][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12685_ (.D(_00564_),
    .CLK(clknet_leaf_193_clock),
    .Q(\u2.mem[35][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12686_ (.D(_00565_),
    .CLK(clknet_leaf_193_clock),
    .Q(\u2.mem[35][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12687_ (.D(_00566_),
    .CLK(clknet_leaf_175_clock),
    .Q(\u2.mem[35][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12688_ (.D(_00567_),
    .CLK(clknet_leaf_177_clock),
    .Q(\u2.mem[35][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12689_ (.D(_00568_),
    .CLK(clknet_leaf_174_clock),
    .Q(\u2.mem[35][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12690_ (.D(_00569_),
    .CLK(clknet_5_27_0_clock),
    .Q(\u2.mem[35][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12691_ (.D(_00570_),
    .CLK(clknet_leaf_89_clock),
    .Q(\u2.mem[35][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12692_ (.D(_00571_),
    .CLK(clknet_leaf_89_clock),
    .Q(\u2.mem[35][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12693_ (.D(_00572_),
    .CLK(clknet_leaf_92_clock),
    .Q(\u2.mem[35][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12694_ (.D(_00573_),
    .CLK(clknet_leaf_92_clock),
    .Q(\u2.mem[35][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12695_ (.D(_00574_),
    .CLK(clknet_leaf_110_clock),
    .Q(\u2.mem[35][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12696_ (.D(_00575_),
    .CLK(clknet_leaf_129_clock),
    .Q(\u2.mem[35][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12697_ (.D(_00576_),
    .CLK(clknet_leaf_111_clock),
    .Q(\u2.mem[35][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12698_ (.D(_00577_),
    .CLK(clknet_leaf_110_clock),
    .Q(\u2.mem[35][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12699_ (.D(_00578_),
    .CLK(clknet_leaf_255_clock),
    .Q(\u2.mem[36][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12700_ (.D(_00579_),
    .CLK(clknet_leaf_256_clock),
    .Q(\u2.mem[36][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12701_ (.D(_00580_),
    .CLK(clknet_leaf_257_clock),
    .Q(\u2.mem[36][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12702_ (.D(_00581_),
    .CLK(clknet_leaf_256_clock),
    .Q(\u2.mem[36][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12703_ (.D(_00582_),
    .CLK(clknet_leaf_239_clock),
    .Q(\u2.mem[36][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12704_ (.D(_00583_),
    .CLK(clknet_leaf_238_clock),
    .Q(\u2.mem[36][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12705_ (.D(_00584_),
    .CLK(clknet_leaf_238_clock),
    .Q(\u2.mem[36][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12706_ (.D(_00585_),
    .CLK(clknet_leaf_238_clock),
    .Q(\u2.mem[36][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12707_ (.D(_00586_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u2.mem[36][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12708_ (.D(_00587_),
    .CLK(clknet_leaf_68_clock),
    .Q(\u2.mem[36][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12709_ (.D(_00588_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u2.mem[36][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12710_ (.D(_00589_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u2.mem[36][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12711_ (.D(_00590_),
    .CLK(clknet_leaf_48_clock),
    .Q(\u2.mem[36][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12712_ (.D(_00591_),
    .CLK(clknet_leaf_50_clock),
    .Q(\u2.mem[36][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12713_ (.D(_00592_),
    .CLK(clknet_leaf_50_clock),
    .Q(\u2.mem[36][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12714_ (.D(_00593_),
    .CLK(clknet_leaf_49_clock),
    .Q(\u2.mem[36][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12715_ (.D(_00594_),
    .CLK(clknet_leaf_252_clock),
    .Q(\u2.mem[37][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12716_ (.D(_00595_),
    .CLK(clknet_leaf_254_clock),
    .Q(\u2.mem[37][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12717_ (.D(_00596_),
    .CLK(clknet_leaf_254_clock),
    .Q(\u2.mem[37][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12718_ (.D(_00597_),
    .CLK(clknet_leaf_252_clock),
    .Q(\u2.mem[37][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12719_ (.D(_00598_),
    .CLK(clknet_leaf_236_clock),
    .Q(\u2.mem[37][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12720_ (.D(_00599_),
    .CLK(clknet_leaf_236_clock),
    .Q(\u2.mem[37][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12721_ (.D(_00600_),
    .CLK(clknet_leaf_235_clock),
    .Q(\u2.mem[37][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12722_ (.D(_00601_),
    .CLK(clknet_leaf_235_clock),
    .Q(\u2.mem[37][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12723_ (.D(_00602_),
    .CLK(clknet_leaf_71_clock),
    .Q(\u2.mem[37][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12724_ (.D(_00603_),
    .CLK(clknet_leaf_72_clock),
    .Q(\u2.mem[37][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12725_ (.D(_00604_),
    .CLK(clknet_leaf_72_clock),
    .Q(\u2.mem[37][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12726_ (.D(_00605_),
    .CLK(clknet_leaf_72_clock),
    .Q(\u2.mem[37][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12727_ (.D(_00606_),
    .CLK(clknet_leaf_43_clock),
    .Q(\u2.mem[37][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12728_ (.D(_00607_),
    .CLK(clknet_leaf_54_clock),
    .Q(\u2.mem[37][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12729_ (.D(_00608_),
    .CLK(clknet_leaf_44_clock),
    .Q(\u2.mem[37][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12730_ (.D(_00609_),
    .CLK(clknet_leaf_43_clock),
    .Q(\u2.mem[37][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12731_ (.D(_00610_),
    .CLK(clknet_leaf_216_clock),
    .Q(\u2.mem[38][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12732_ (.D(_00611_),
    .CLK(clknet_leaf_255_clock),
    .Q(\u2.mem[38][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12733_ (.D(_00612_),
    .CLK(clknet_leaf_255_clock),
    .Q(\u2.mem[38][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12734_ (.D(_00613_),
    .CLK(clknet_leaf_252_clock),
    .Q(\u2.mem[38][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12735_ (.D(_00614_),
    .CLK(clknet_leaf_237_clock),
    .Q(\u2.mem[38][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12736_ (.D(_00615_),
    .CLK(clknet_leaf_229_clock),
    .Q(\u2.mem[38][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12737_ (.D(_00616_),
    .CLK(clknet_leaf_232_clock),
    .Q(\u2.mem[38][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12738_ (.D(_00617_),
    .CLK(clknet_leaf_234_clock),
    .Q(\u2.mem[38][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12739_ (.D(_00618_),
    .CLK(clknet_leaf_65_clock),
    .Q(\u2.mem[38][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12740_ (.D(_00619_),
    .CLK(clknet_leaf_67_clock),
    .Q(\u2.mem[38][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12741_ (.D(_00620_),
    .CLK(clknet_leaf_70_clock),
    .Q(\u2.mem[38][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12742_ (.D(_00621_),
    .CLK(clknet_leaf_70_clock),
    .Q(\u2.mem[38][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12743_ (.D(_00622_),
    .CLK(clknet_leaf_53_clock),
    .Q(\u2.mem[38][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12744_ (.D(_00623_),
    .CLK(clknet_leaf_50_clock),
    .Q(\u2.mem[38][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12745_ (.D(_00624_),
    .CLK(clknet_leaf_53_clock),
    .Q(\u2.mem[38][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12746_ (.D(_00625_),
    .CLK(clknet_leaf_50_clock),
    .Q(\u2.mem[38][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12747_ (.D(_00626_),
    .CLK(clknet_leaf_216_clock),
    .Q(\u2.mem[39][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12748_ (.D(_00627_),
    .CLK(clknet_leaf_211_clock),
    .Q(\u2.mem[39][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12749_ (.D(_00628_),
    .CLK(clknet_leaf_212_clock),
    .Q(\u2.mem[39][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12750_ (.D(_00629_),
    .CLK(clknet_leaf_213_clock),
    .Q(\u2.mem[39][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12751_ (.D(_00630_),
    .CLK(clknet_leaf_225_clock),
    .Q(\u2.mem[39][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12752_ (.D(_00631_),
    .CLK(clknet_leaf_227_clock),
    .Q(\u2.mem[39][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12753_ (.D(_00632_),
    .CLK(clknet_leaf_230_clock),
    .Q(\u2.mem[39][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12754_ (.D(_00633_),
    .CLK(clknet_leaf_229_clock),
    .Q(\u2.mem[39][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12755_ (.D(_00634_),
    .CLK(clknet_leaf_64_clock),
    .Q(\u2.mem[39][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12756_ (.D(_00635_),
    .CLK(clknet_leaf_69_clock),
    .Q(\u2.mem[39][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12757_ (.D(_00636_),
    .CLK(clknet_leaf_70_clock),
    .Q(\u2.mem[39][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12758_ (.D(_00637_),
    .CLK(clknet_leaf_74_clock),
    .Q(\u2.mem[39][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12759_ (.D(_00638_),
    .CLK(clknet_leaf_50_clock),
    .Q(\u2.mem[39][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12760_ (.D(_00639_),
    .CLK(clknet_leaf_51_clock),
    .Q(\u2.mem[39][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12761_ (.D(_00640_),
    .CLK(clknet_leaf_141_clock),
    .Q(\u2.mem[39][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12762_ (.D(_00641_),
    .CLK(clknet_5_13_0_clock),
    .Q(\u2.mem[39][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12763_ (.D(_00642_),
    .CLK(clknet_leaf_203_clock),
    .Q(\u2.mem[40][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12764_ (.D(_00643_),
    .CLK(clknet_leaf_203_clock),
    .Q(\u2.mem[40][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12765_ (.D(_00644_),
    .CLK(clknet_leaf_204_clock),
    .Q(\u2.mem[40][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12766_ (.D(_00645_),
    .CLK(clknet_leaf_203_clock),
    .Q(\u2.mem[40][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12767_ (.D(_00646_),
    .CLK(clknet_leaf_155_clock),
    .Q(\u2.mem[40][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12768_ (.D(_00647_),
    .CLK(clknet_leaf_155_clock),
    .Q(\u2.mem[40][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12769_ (.D(_00648_),
    .CLK(clknet_leaf_154_clock),
    .Q(\u2.mem[40][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12770_ (.D(_00649_),
    .CLK(clknet_leaf_155_clock),
    .Q(\u2.mem[40][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12771_ (.D(_00650_),
    .CLK(clknet_leaf_90_clock),
    .Q(\u2.mem[40][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12772_ (.D(_00651_),
    .CLK(clknet_leaf_91_clock),
    .Q(\u2.mem[40][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12773_ (.D(_00652_),
    .CLK(clknet_leaf_79_clock),
    .Q(\u2.mem[40][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12774_ (.D(_00653_),
    .CLK(clknet_leaf_79_clock),
    .Q(\u2.mem[40][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12775_ (.D(_00654_),
    .CLK(clknet_leaf_131_clock),
    .Q(\u2.mem[40][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12776_ (.D(_00655_),
    .CLK(clknet_leaf_130_clock),
    .Q(\u2.mem[40][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12777_ (.D(_00656_),
    .CLK(clknet_leaf_130_clock),
    .Q(\u2.mem[40][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12778_ (.D(_00657_),
    .CLK(clknet_leaf_130_clock),
    .Q(\u2.mem[40][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12779_ (.D(_00658_),
    .CLK(clknet_leaf_253_clock),
    .Q(\u2.mem[41][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12780_ (.D(_00659_),
    .CLK(clknet_leaf_253_clock),
    .Q(\u2.mem[41][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12781_ (.D(_00660_),
    .CLK(clknet_leaf_253_clock),
    .Q(\u2.mem[41][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12782_ (.D(_00661_),
    .CLK(clknet_leaf_253_clock),
    .Q(\u2.mem[41][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12783_ (.D(_00662_),
    .CLK(clknet_leaf_322_clock),
    .Q(\u2.mem[41][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12784_ (.D(_00663_),
    .CLK(clknet_leaf_321_clock),
    .Q(\u2.mem[41][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12785_ (.D(_00664_),
    .CLK(clknet_leaf_235_clock),
    .Q(\u2.mem[41][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12786_ (.D(_00665_),
    .CLK(clknet_leaf_321_clock),
    .Q(\u2.mem[41][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12787_ (.D(_00666_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u2.mem[41][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12788_ (.D(_00667_),
    .CLK(clknet_leaf_71_clock),
    .Q(\u2.mem[41][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12789_ (.D(_00668_),
    .CLK(clknet_leaf_71_clock),
    .Q(\u2.mem[41][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12790_ (.D(_00669_),
    .CLK(clknet_leaf_71_clock),
    .Q(\u2.mem[41][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12791_ (.D(_00670_),
    .CLK(clknet_leaf_44_clock),
    .Q(\u2.mem[41][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12792_ (.D(_00671_),
    .CLK(clknet_leaf_44_clock),
    .Q(\u2.mem[41][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12793_ (.D(_00672_),
    .CLK(clknet_leaf_48_clock),
    .Q(\u2.mem[41][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12794_ (.D(_00673_),
    .CLK(clknet_leaf_48_clock),
    .Q(\u2.mem[41][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12795_ (.D(_00674_),
    .CLK(clknet_leaf_220_clock),
    .Q(\u2.mem[42][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12796_ (.D(_00675_),
    .CLK(clknet_leaf_220_clock),
    .Q(\u2.mem[42][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12797_ (.D(_00676_),
    .CLK(clknet_leaf_220_clock),
    .Q(\u2.mem[42][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12798_ (.D(_00677_),
    .CLK(clknet_leaf_220_clock),
    .Q(\u2.mem[42][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12799_ (.D(_00678_),
    .CLK(clknet_leaf_144_clock),
    .Q(\u2.mem[42][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12800_ (.D(_00679_),
    .CLK(clknet_leaf_144_clock),
    .Q(\u2.mem[42][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12801_ (.D(_00680_),
    .CLK(clknet_leaf_144_clock),
    .Q(\u2.mem[42][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12802_ (.D(_00681_),
    .CLK(clknet_leaf_145_clock),
    .Q(\u2.mem[42][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12803_ (.D(_00682_),
    .CLK(clknet_leaf_145_clock),
    .Q(\u2.mem[42][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12804_ (.D(_00683_),
    .CLK(clknet_leaf_62_clock),
    .Q(\u2.mem[42][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12805_ (.D(_00684_),
    .CLK(clknet_leaf_82_clock),
    .Q(\u2.mem[42][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12806_ (.D(_00685_),
    .CLK(clknet_leaf_82_clock),
    .Q(\u2.mem[42][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12807_ (.D(_00686_),
    .CLK(clknet_leaf_140_clock),
    .Q(\u2.mem[42][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12808_ (.D(_00687_),
    .CLK(clknet_leaf_139_clock),
    .Q(\u2.mem[42][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12809_ (.D(_00688_),
    .CLK(clknet_leaf_139_clock),
    .Q(\u2.mem[42][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12810_ (.D(_00689_),
    .CLK(clknet_leaf_139_clock),
    .Q(\u2.mem[42][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12811_ (.D(_00690_),
    .CLK(clknet_leaf_221_clock),
    .Q(\u2.mem[43][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12812_ (.D(_00691_),
    .CLK(clknet_leaf_201_clock),
    .Q(\u2.mem[43][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12813_ (.D(_00692_),
    .CLK(clknet_leaf_201_clock),
    .Q(\u2.mem[43][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12814_ (.D(_00693_),
    .CLK(clknet_leaf_220_clock),
    .Q(\u2.mem[43][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12815_ (.D(_00694_),
    .CLK(clknet_leaf_146_clock),
    .Q(\u2.mem[43][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12816_ (.D(_00695_),
    .CLK(clknet_leaf_147_clock),
    .Q(\u2.mem[43][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12817_ (.D(_00696_),
    .CLK(clknet_leaf_146_clock),
    .Q(\u2.mem[43][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12818_ (.D(_00697_),
    .CLK(clknet_leaf_147_clock),
    .Q(\u2.mem[43][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12819_ (.D(_00698_),
    .CLK(clknet_leaf_60_clock),
    .Q(\u2.mem[43][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12820_ (.D(_00699_),
    .CLK(clknet_leaf_61_clock),
    .Q(\u2.mem[43][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12821_ (.D(_00700_),
    .CLK(clknet_leaf_83_clock),
    .Q(\u2.mem[43][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12822_ (.D(_00701_),
    .CLK(clknet_leaf_83_clock),
    .Q(\u2.mem[43][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12823_ (.D(_00702_),
    .CLK(clknet_leaf_135_clock),
    .Q(\u2.mem[43][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12824_ (.D(_00703_),
    .CLK(clknet_leaf_137_clock),
    .Q(\u2.mem[43][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12825_ (.D(_00704_),
    .CLK(clknet_leaf_136_clock),
    .Q(\u2.mem[43][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12826_ (.D(_00705_),
    .CLK(clknet_leaf_136_clock),
    .Q(\u2.mem[43][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12827_ (.D(_00706_),
    .CLK(clknet_leaf_221_clock),
    .Q(\u2.mem[44][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12828_ (.D(_00707_),
    .CLK(clknet_leaf_208_clock),
    .Q(\u2.mem[44][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12829_ (.D(_00708_),
    .CLK(clknet_leaf_207_clock),
    .Q(\u2.mem[44][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12830_ (.D(_00709_),
    .CLK(clknet_leaf_220_clock),
    .Q(\u2.mem[44][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12831_ (.D(_00710_),
    .CLK(clknet_leaf_149_clock),
    .Q(\u2.mem[44][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12832_ (.D(_00711_),
    .CLK(clknet_leaf_145_clock),
    .Q(\u2.mem[44][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12833_ (.D(_00712_),
    .CLK(clknet_leaf_148_clock),
    .Q(\u2.mem[44][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12834_ (.D(_00713_),
    .CLK(clknet_leaf_145_clock),
    .Q(\u2.mem[44][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12835_ (.D(_00714_),
    .CLK(clknet_leaf_146_clock),
    .Q(\u2.mem[44][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12836_ (.D(_00715_),
    .CLK(clknet_leaf_61_clock),
    .Q(\u2.mem[44][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12837_ (.D(_00716_),
    .CLK(clknet_leaf_82_clock),
    .Q(\u2.mem[44][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12838_ (.D(_00717_),
    .CLK(clknet_leaf_63_clock),
    .Q(\u2.mem[44][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12839_ (.D(_00718_),
    .CLK(clknet_leaf_135_clock),
    .Q(\u2.mem[44][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12840_ (.D(_00719_),
    .CLK(clknet_leaf_139_clock),
    .Q(\u2.mem[44][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12841_ (.D(_00720_),
    .CLK(clknet_leaf_138_clock),
    .Q(\u2.mem[44][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12842_ (.D(_00721_),
    .CLK(clknet_leaf_139_clock),
    .Q(\u2.mem[44][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12843_ (.D(_00722_),
    .CLK(clknet_leaf_198_clock),
    .Q(\u2.mem[45][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12844_ (.D(_00723_),
    .CLK(clknet_leaf_204_clock),
    .Q(\u2.mem[45][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12845_ (.D(_00724_),
    .CLK(clknet_leaf_205_clock),
    .Q(\u2.mem[45][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12846_ (.D(_00725_),
    .CLK(clknet_leaf_203_clock),
    .Q(\u2.mem[45][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12847_ (.D(_00726_),
    .CLK(clknet_leaf_151_clock),
    .Q(\u2.mem[45][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12848_ (.D(_00727_),
    .CLK(clknet_leaf_151_clock),
    .Q(\u2.mem[45][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12849_ (.D(_00728_),
    .CLK(clknet_leaf_154_clock),
    .Q(\u2.mem[45][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12850_ (.D(_00729_),
    .CLK(clknet_leaf_150_clock),
    .Q(\u2.mem[45][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12851_ (.D(_00730_),
    .CLK(clknet_leaf_86_clock),
    .Q(\u2.mem[45][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12852_ (.D(_00731_),
    .CLK(clknet_leaf_90_clock),
    .Q(\u2.mem[45][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12853_ (.D(_00732_),
    .CLK(clknet_leaf_80_clock),
    .Q(\u2.mem[45][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12854_ (.D(_00733_),
    .CLK(clknet_leaf_80_clock),
    .Q(\u2.mem[45][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12855_ (.D(_00734_),
    .CLK(clknet_leaf_133_clock),
    .Q(\u2.mem[45][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12856_ (.D(_00735_),
    .CLK(clknet_leaf_129_clock),
    .Q(\u2.mem[45][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12857_ (.D(_00736_),
    .CLK(clknet_leaf_133_clock),
    .Q(\u2.mem[45][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12858_ (.D(_00737_),
    .CLK(clknet_leaf_129_clock),
    .Q(\u2.mem[45][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12859_ (.D(_00738_),
    .CLK(clknet_leaf_199_clock),
    .Q(\u2.mem[46][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12860_ (.D(_00739_),
    .CLK(clknet_leaf_203_clock),
    .Q(\u2.mem[46][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12861_ (.D(_00740_),
    .CLK(clknet_leaf_200_clock),
    .Q(\u2.mem[46][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12862_ (.D(_00741_),
    .CLK(clknet_leaf_199_clock),
    .Q(\u2.mem[46][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12863_ (.D(_00742_),
    .CLK(clknet_leaf_148_clock),
    .Q(\u2.mem[46][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12864_ (.D(_00743_),
    .CLK(clknet_leaf_148_clock),
    .Q(\u2.mem[46][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12865_ (.D(_00744_),
    .CLK(clknet_leaf_148_clock),
    .Q(\u2.mem[46][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12866_ (.D(_00745_),
    .CLK(clknet_leaf_151_clock),
    .Q(\u2.mem[46][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12867_ (.D(_00746_),
    .CLK(clknet_leaf_60_clock),
    .Q(\u2.mem[46][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12868_ (.D(_00747_),
    .CLK(clknet_leaf_83_clock),
    .Q(\u2.mem[46][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12869_ (.D(_00748_),
    .CLK(clknet_leaf_80_clock),
    .Q(\u2.mem[46][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12870_ (.D(_00749_),
    .CLK(clknet_leaf_83_clock),
    .Q(\u2.mem[46][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12871_ (.D(_00750_),
    .CLK(clknet_leaf_136_clock),
    .Q(\u2.mem[46][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12872_ (.D(_00751_),
    .CLK(clknet_leaf_137_clock),
    .Q(\u2.mem[46][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12873_ (.D(_00752_),
    .CLK(clknet_leaf_137_clock),
    .Q(\u2.mem[46][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12874_ (.D(_00753_),
    .CLK(clknet_leaf_137_clock),
    .Q(\u2.mem[46][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12875_ (.D(_00754_),
    .CLK(clknet_leaf_218_clock),
    .Q(\u2.mem[47][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12876_ (.D(_00755_),
    .CLK(clknet_leaf_215_clock),
    .Q(\u2.mem[47][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12877_ (.D(_00756_),
    .CLK(clknet_leaf_214_clock),
    .Q(\u2.mem[47][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12878_ (.D(_00757_),
    .CLK(clknet_leaf_219_clock),
    .Q(\u2.mem[47][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12879_ (.D(_00758_),
    .CLK(clknet_leaf_230_clock),
    .Q(\u2.mem[47][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12880_ (.D(_00759_),
    .CLK(clknet_leaf_230_clock),
    .Q(\u2.mem[47][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12881_ (.D(_00760_),
    .CLK(clknet_leaf_143_clock),
    .Q(\u2.mem[47][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12882_ (.D(_00761_),
    .CLK(clknet_leaf_230_clock),
    .Q(\u2.mem[47][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12883_ (.D(_00762_),
    .CLK(clknet_leaf_64_clock),
    .Q(\u2.mem[47][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12884_ (.D(_00763_),
    .CLK(clknet_leaf_63_clock),
    .Q(\u2.mem[47][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12885_ (.D(_00764_),
    .CLK(clknet_leaf_63_clock),
    .Q(\u2.mem[47][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12886_ (.D(_00765_),
    .CLK(clknet_leaf_63_clock),
    .Q(\u2.mem[47][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12887_ (.D(_00766_),
    .CLK(clknet_leaf_57_clock),
    .Q(\u2.mem[47][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12888_ (.D(_00767_),
    .CLK(clknet_leaf_57_clock),
    .Q(\u2.mem[47][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12889_ (.D(_00768_),
    .CLK(clknet_leaf_51_clock),
    .Q(\u2.mem[47][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12890_ (.D(_00769_),
    .CLK(clknet_leaf_140_clock),
    .Q(\u2.mem[47][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12891_ (.D(_00770_),
    .CLK(clknet_leaf_219_clock),
    .Q(\u2.mem[48][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12892_ (.D(_00771_),
    .CLK(clknet_leaf_209_clock),
    .Q(\u2.mem[48][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12893_ (.D(_00772_),
    .CLK(clknet_leaf_214_clock),
    .Q(\u2.mem[48][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12894_ (.D(_00773_),
    .CLK(clknet_leaf_214_clock),
    .Q(\u2.mem[48][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12895_ (.D(_00774_),
    .CLK(clknet_leaf_225_clock),
    .Q(\u2.mem[48][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12896_ (.D(_00775_),
    .CLK(clknet_leaf_224_clock),
    .Q(\u2.mem[48][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12897_ (.D(_00776_),
    .CLK(clknet_leaf_224_clock),
    .Q(\u2.mem[48][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12898_ (.D(_00777_),
    .CLK(clknet_leaf_230_clock),
    .Q(\u2.mem[48][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12899_ (.D(_00778_),
    .CLK(clknet_leaf_64_clock),
    .Q(\u2.mem[48][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12900_ (.D(_00779_),
    .CLK(clknet_leaf_75_clock),
    .Q(\u2.mem[48][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12901_ (.D(_00780_),
    .CLK(clknet_leaf_74_clock),
    .Q(\u2.mem[48][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12902_ (.D(_00781_),
    .CLK(clknet_leaf_74_clock),
    .Q(\u2.mem[48][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12903_ (.D(_00782_),
    .CLK(clknet_leaf_140_clock),
    .Q(\u2.mem[48][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12904_ (.D(_00783_),
    .CLK(clknet_leaf_51_clock),
    .Q(\u2.mem[48][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12905_ (.D(_00784_),
    .CLK(clknet_leaf_141_clock),
    .Q(\u2.mem[48][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12906_ (.D(_00785_),
    .CLK(clknet_leaf_141_clock),
    .Q(\u2.mem[48][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12907_ (.D(_00786_),
    .CLK(clknet_leaf_221_clock),
    .Q(\u2.mem[49][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12908_ (.D(_00787_),
    .CLK(clknet_leaf_202_clock),
    .Q(\u2.mem[49][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12909_ (.D(_00788_),
    .CLK(clknet_leaf_202_clock),
    .Q(\u2.mem[49][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12910_ (.D(_00789_),
    .CLK(clknet_leaf_202_clock),
    .Q(\u2.mem[49][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12911_ (.D(_00790_),
    .CLK(clknet_leaf_157_clock),
    .Q(\u2.mem[49][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12912_ (.D(_00791_),
    .CLK(clknet_leaf_147_clock),
    .Q(\u2.mem[49][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12913_ (.D(_00792_),
    .CLK(clknet_leaf_158_clock),
    .Q(\u2.mem[49][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12914_ (.D(_00793_),
    .CLK(clknet_leaf_157_clock),
    .Q(\u2.mem[49][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12915_ (.D(_00794_),
    .CLK(clknet_leaf_147_clock),
    .Q(\u2.mem[49][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12916_ (.D(_00795_),
    .CLK(clknet_leaf_60_clock),
    .Q(\u2.mem[49][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12917_ (.D(_00796_),
    .CLK(clknet_leaf_83_clock),
    .Q(\u2.mem[49][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12918_ (.D(_00797_),
    .CLK(clknet_leaf_84_clock),
    .Q(\u2.mem[49][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12919_ (.D(_00798_),
    .CLK(clknet_leaf_125_clock),
    .Q(\u2.mem[49][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12920_ (.D(_00799_),
    .CLK(clknet_leaf_138_clock),
    .Q(\u2.mem[49][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12921_ (.D(_00800_),
    .CLK(clknet_leaf_159_clock),
    .Q(\u2.mem[49][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12922_ (.D(_00801_),
    .CLK(clknet_leaf_126_clock),
    .Q(\u2.mem[49][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12923_ (.D(_00802_),
    .CLK(clknet_leaf_252_clock),
    .Q(\u2.mem[50][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12924_ (.D(_00803_),
    .CLK(clknet_leaf_257_clock),
    .Q(\u2.mem[50][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12925_ (.D(_00804_),
    .CLK(clknet_leaf_257_clock),
    .Q(\u2.mem[50][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12926_ (.D(_00805_),
    .CLK(clknet_leaf_255_clock),
    .Q(\u2.mem[50][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12927_ (.D(_00806_),
    .CLK(clknet_leaf_234_clock),
    .Q(\u2.mem[50][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12928_ (.D(_00807_),
    .CLK(clknet_leaf_235_clock),
    .Q(\u2.mem[50][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12929_ (.D(_00808_),
    .CLK(clknet_leaf_233_clock),
    .Q(\u2.mem[50][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12930_ (.D(_00809_),
    .CLK(clknet_leaf_234_clock),
    .Q(\u2.mem[50][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12931_ (.D(_00810_),
    .CLK(clknet_leaf_232_clock),
    .Q(\u2.mem[50][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12932_ (.D(_00811_),
    .CLK(clknet_leaf_66_clock),
    .Q(\u2.mem[50][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12933_ (.D(_00812_),
    .CLK(clknet_leaf_67_clock),
    .Q(\u2.mem[50][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12934_ (.D(_00813_),
    .CLK(clknet_leaf_31_clock),
    .Q(\u2.mem[50][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12935_ (.D(_00814_),
    .CLK(clknet_leaf_49_clock),
    .Q(\u2.mem[50][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12936_ (.D(_00815_),
    .CLK(clknet_leaf_324_clock),
    .Q(\u2.mem[50][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12937_ (.D(_00816_),
    .CLK(clknet_leaf_323_clock),
    .Q(\u2.mem[50][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12938_ (.D(_00817_),
    .CLK(clknet_leaf_325_clock),
    .Q(\u2.mem[50][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12939_ (.D(_00818_),
    .CLK(clknet_leaf_251_clock),
    .Q(\u2.mem[51][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12940_ (.D(_00819_),
    .CLK(clknet_leaf_256_clock),
    .Q(\u2.mem[51][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12941_ (.D(_00820_),
    .CLK(clknet_leaf_256_clock),
    .Q(\u2.mem[51][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12942_ (.D(_00821_),
    .CLK(clknet_leaf_255_clock),
    .Q(\u2.mem[51][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12943_ (.D(_00822_),
    .CLK(clknet_leaf_237_clock),
    .Q(\u2.mem[51][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12944_ (.D(_00823_),
    .CLK(clknet_leaf_235_clock),
    .Q(\u2.mem[51][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12945_ (.D(_00824_),
    .CLK(clknet_leaf_233_clock),
    .Q(\u2.mem[51][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12946_ (.D(_00825_),
    .CLK(clknet_leaf_233_clock),
    .Q(\u2.mem[51][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12947_ (.D(_00826_),
    .CLK(clknet_leaf_233_clock),
    .Q(\u2.mem[51][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12948_ (.D(_00827_),
    .CLK(clknet_leaf_66_clock),
    .Q(\u2.mem[51][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12949_ (.D(_00828_),
    .CLK(clknet_leaf_67_clock),
    .Q(\u2.mem[51][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12950_ (.D(_00829_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u2.mem[51][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12951_ (.D(_00830_),
    .CLK(clknet_leaf_49_clock),
    .Q(\u2.mem[51][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12952_ (.D(_00831_),
    .CLK(clknet_leaf_49_clock),
    .Q(\u2.mem[51][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12953_ (.D(_00832_),
    .CLK(clknet_leaf_324_clock),
    .Q(\u2.mem[51][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12954_ (.D(_00833_),
    .CLK(clknet_leaf_324_clock),
    .Q(\u2.mem[51][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12955_ (.D(_00834_),
    .CLK(clknet_leaf_198_clock),
    .Q(\u2.mem[52][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12956_ (.D(_00835_),
    .CLK(clknet_leaf_197_clock),
    .Q(\u2.mem[52][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12957_ (.D(_00836_),
    .CLK(clknet_leaf_196_clock),
    .Q(\u2.mem[52][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12958_ (.D(_00837_),
    .CLK(clknet_leaf_197_clock),
    .Q(\u2.mem[52][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12959_ (.D(_00838_),
    .CLK(clknet_leaf_155_clock),
    .Q(\u2.mem[52][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12960_ (.D(_00839_),
    .CLK(clknet_leaf_156_clock),
    .Q(\u2.mem[52][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12961_ (.D(_00840_),
    .CLK(clknet_leaf_157_clock),
    .Q(\u2.mem[52][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12962_ (.D(_00841_),
    .CLK(clknet_leaf_156_clock),
    .Q(\u2.mem[52][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12963_ (.D(_00842_),
    .CLK(clknet_leaf_109_clock),
    .Q(\u2.mem[52][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12964_ (.D(_00843_),
    .CLK(clknet_leaf_109_clock),
    .Q(\u2.mem[52][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12965_ (.D(_00844_),
    .CLK(clknet_leaf_85_clock),
    .Q(\u2.mem[52][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12966_ (.D(_00845_),
    .CLK(clknet_leaf_87_clock),
    .Q(\u2.mem[52][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12967_ (.D(_00846_),
    .CLK(clknet_leaf_124_clock),
    .Q(\u2.mem[52][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12968_ (.D(_00847_),
    .CLK(clknet_leaf_124_clock),
    .Q(\u2.mem[52][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12969_ (.D(_00848_),
    .CLK(clknet_leaf_125_clock),
    .Q(\u2.mem[52][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12970_ (.D(_00849_),
    .CLK(clknet_leaf_124_clock),
    .Q(\u2.mem[52][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12971_ (.D(_00850_),
    .CLK(clknet_leaf_246_clock),
    .Q(\u2.mem[53][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12972_ (.D(_00851_),
    .CLK(clknet_leaf_262_clock),
    .Q(\u2.mem[53][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12973_ (.D(_00852_),
    .CLK(clknet_leaf_262_clock),
    .Q(\u2.mem[53][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12974_ (.D(_00853_),
    .CLK(clknet_leaf_261_clock),
    .Q(\u2.mem[53][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12975_ (.D(_00854_),
    .CLK(clknet_leaf_249_clock),
    .Q(\u2.mem[53][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12976_ (.D(_00855_),
    .CLK(clknet_leaf_249_clock),
    .Q(\u2.mem[53][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12977_ (.D(_00856_),
    .CLK(clknet_leaf_250_clock),
    .Q(\u2.mem[53][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12978_ (.D(_00857_),
    .CLK(clknet_leaf_250_clock),
    .Q(\u2.mem[53][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12979_ (.D(_00858_),
    .CLK(clknet_leaf_42_clock),
    .Q(\u2.mem[53][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12980_ (.D(_00859_),
    .CLK(clknet_leaf_43_clock),
    .Q(\u2.mem[53][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12981_ (.D(_00860_),
    .CLK(clknet_leaf_31_clock),
    .Q(\u2.mem[53][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12982_ (.D(_00861_),
    .CLK(clknet_leaf_31_clock),
    .Q(\u2.mem[53][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12983_ (.D(_00862_),
    .CLK(clknet_leaf_326_clock),
    .Q(\u2.mem[53][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12984_ (.D(_00863_),
    .CLK(clknet_leaf_329_clock),
    .Q(\u2.mem[53][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12985_ (.D(_00864_),
    .CLK(clknet_leaf_319_clock),
    .Q(\u2.mem[53][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12986_ (.D(_00865_),
    .CLK(clknet_leaf_326_clock),
    .Q(\u2.mem[53][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12987_ (.D(_00866_),
    .CLK(clknet_leaf_248_clock),
    .Q(\u2.mem[54][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12988_ (.D(_00867_),
    .CLK(clknet_leaf_257_clock),
    .Q(\u2.mem[54][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12989_ (.D(_00868_),
    .CLK(clknet_leaf_258_clock),
    .Q(\u2.mem[54][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12990_ (.D(_00869_),
    .CLK(clknet_leaf_258_clock),
    .Q(\u2.mem[54][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12991_ (.D(_00870_),
    .CLK(clknet_leaf_239_clock),
    .Q(\u2.mem[54][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12992_ (.D(_00871_),
    .CLK(clknet_leaf_240_clock),
    .Q(\u2.mem[54][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12993_ (.D(_00872_),
    .CLK(clknet_leaf_239_clock),
    .Q(\u2.mem[54][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12994_ (.D(_00873_),
    .CLK(clknet_leaf_236_clock),
    .Q(\u2.mem[54][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12995_ (.D(_00874_),
    .CLK(clknet_leaf_323_clock),
    .Q(\u2.mem[54][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12996_ (.D(_00875_),
    .CLK(clknet_leaf_33_clock),
    .Q(\u2.mem[54][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12997_ (.D(_00876_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u2.mem[54][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12998_ (.D(_00877_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u2.mem[54][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12999_ (.D(_00878_),
    .CLK(clknet_leaf_323_clock),
    .Q(\u2.mem[54][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13000_ (.D(_00879_),
    .CLK(clknet_leaf_322_clock),
    .Q(\u2.mem[54][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13001_ (.D(_00880_),
    .CLK(clknet_leaf_322_clock),
    .Q(\u2.mem[54][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13002_ (.D(_00881_),
    .CLK(clknet_leaf_322_clock),
    .Q(\u2.mem[54][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13003_ (.D(_00882_),
    .CLK(clknet_leaf_249_clock),
    .Q(\u2.mem[55][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13004_ (.D(_00883_),
    .CLK(clknet_leaf_257_clock),
    .Q(\u2.mem[55][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13005_ (.D(_00884_),
    .CLK(clknet_leaf_258_clock),
    .Q(\u2.mem[55][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13006_ (.D(_00885_),
    .CLK(clknet_leaf_259_clock),
    .Q(\u2.mem[55][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13007_ (.D(_00886_),
    .CLK(clknet_leaf_240_clock),
    .Q(\u2.mem[55][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13008_ (.D(_00887_),
    .CLK(clknet_leaf_240_clock),
    .Q(\u2.mem[55][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13009_ (.D(_00888_),
    .CLK(clknet_leaf_239_clock),
    .Q(\u2.mem[55][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13010_ (.D(_00889_),
    .CLK(clknet_leaf_237_clock),
    .Q(\u2.mem[55][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13011_ (.D(_00890_),
    .CLK(clknet_leaf_323_clock),
    .Q(\u2.mem[55][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13012_ (.D(_00891_),
    .CLK(clknet_leaf_31_clock),
    .Q(\u2.mem[55][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13013_ (.D(_00892_),
    .CLK(clknet_leaf_29_clock),
    .Q(\u2.mem[55][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13014_ (.D(_00893_),
    .CLK(clknet_leaf_28_clock),
    .Q(\u2.mem[55][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13015_ (.D(_00894_),
    .CLK(clknet_leaf_323_clock),
    .Q(\u2.mem[55][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13016_ (.D(_00895_),
    .CLK(clknet_leaf_319_clock),
    .Q(\u2.mem[55][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13017_ (.D(_00896_),
    .CLK(clknet_leaf_319_clock),
    .Q(\u2.mem[55][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13018_ (.D(_00897_),
    .CLK(clknet_leaf_322_clock),
    .Q(\u2.mem[55][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13019_ (.D(_00898_),
    .CLK(clknet_leaf_249_clock),
    .Q(\u2.mem[56][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13020_ (.D(_00899_),
    .CLK(clknet_leaf_258_clock),
    .Q(\u2.mem[56][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13021_ (.D(_00900_),
    .CLK(clknet_leaf_258_clock),
    .Q(\u2.mem[56][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13022_ (.D(_00901_),
    .CLK(clknet_leaf_259_clock),
    .Q(\u2.mem[56][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13023_ (.D(_00902_),
    .CLK(clknet_leaf_249_clock),
    .Q(\u2.mem[56][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13024_ (.D(_00903_),
    .CLK(clknet_leaf_246_clock),
    .Q(\u2.mem[56][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13025_ (.D(_00904_),
    .CLK(clknet_leaf_251_clock),
    .Q(\u2.mem[56][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13026_ (.D(_00905_),
    .CLK(clknet_leaf_251_clock),
    .Q(\u2.mem[56][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13027_ (.D(_00906_),
    .CLK(clknet_leaf_42_clock),
    .Q(\u2.mem[56][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13028_ (.D(_00907_),
    .CLK(clknet_leaf_31_clock),
    .Q(\u2.mem[56][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13029_ (.D(_00908_),
    .CLK(clknet_leaf_31_clock),
    .Q(\u2.mem[56][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13030_ (.D(_00909_),
    .CLK(clknet_leaf_32_clock),
    .Q(\u2.mem[56][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13031_ (.D(_00910_),
    .CLK(clknet_leaf_326_clock),
    .Q(\u2.mem[56][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13032_ (.D(_00911_),
    .CLK(clknet_leaf_328_clock),
    .Q(\u2.mem[56][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13033_ (.D(_00912_),
    .CLK(clknet_leaf_328_clock),
    .Q(\u2.mem[56][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13034_ (.D(_00913_),
    .CLK(clknet_leaf_326_clock),
    .Q(\u2.mem[56][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13035_ (.D(_00914_),
    .CLK(clknet_leaf_248_clock),
    .Q(\u2.mem[57][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13036_ (.D(_00915_),
    .CLK(clknet_leaf_260_clock),
    .Q(\u2.mem[57][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13037_ (.D(_00916_),
    .CLK(clknet_leaf_267_clock),
    .Q(\u2.mem[57][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13038_ (.D(_00917_),
    .CLK(clknet_leaf_248_clock),
    .Q(\u2.mem[57][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13039_ (.D(_00918_),
    .CLK(clknet_leaf_320_clock),
    .Q(\u2.mem[57][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13040_ (.D(_00919_),
    .CLK(clknet_leaf_320_clock),
    .Q(\u2.mem[57][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13041_ (.D(_00920_),
    .CLK(clknet_leaf_321_clock),
    .Q(\u2.mem[57][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13042_ (.D(_00921_),
    .CLK(clknet_leaf_321_clock),
    .Q(\u2.mem[57][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13043_ (.D(_00922_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u2.mem[57][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13044_ (.D(_00923_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u2.mem[57][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13045_ (.D(_00924_),
    .CLK(clknet_leaf_25_clock),
    .Q(\u2.mem[57][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13046_ (.D(_00925_),
    .CLK(clknet_leaf_25_clock),
    .Q(\u2.mem[57][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13047_ (.D(_00926_),
    .CLK(clknet_leaf_44_clock),
    .Q(\u2.mem[57][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13048_ (.D(_00927_),
    .CLK(clknet_leaf_44_clock),
    .Q(\u2.mem[57][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13049_ (.D(_00928_),
    .CLK(clknet_leaf_45_clock),
    .Q(\u2.mem[57][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13050_ (.D(_00929_),
    .CLK(clknet_leaf_44_clock),
    .Q(\u2.mem[57][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13051_ (.D(_00930_),
    .CLK(clknet_leaf_254_clock),
    .Q(\u2.mem[58][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13052_ (.D(_00931_),
    .CLK(clknet_leaf_259_clock),
    .Q(\u2.mem[58][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13053_ (.D(_00932_),
    .CLK(clknet_leaf_259_clock),
    .Q(\u2.mem[58][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13054_ (.D(_00933_),
    .CLK(clknet_leaf_259_clock),
    .Q(\u2.mem[58][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13055_ (.D(_00934_),
    .CLK(clknet_leaf_240_clock),
    .Q(\u2.mem[58][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13056_ (.D(_00935_),
    .CLK(clknet_leaf_243_clock),
    .Q(\u2.mem[58][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13057_ (.D(_00936_),
    .CLK(clknet_leaf_240_clock),
    .Q(\u2.mem[58][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13058_ (.D(_00937_),
    .CLK(clknet_leaf_242_clock),
    .Q(\u2.mem[58][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13059_ (.D(_00938_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u2.mem[58][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13060_ (.D(_00939_),
    .CLK(clknet_leaf_27_clock),
    .Q(\u2.mem[58][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13061_ (.D(_00940_),
    .CLK(clknet_leaf_26_clock),
    .Q(\u2.mem[58][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13062_ (.D(_00941_),
    .CLK(clknet_leaf_30_clock),
    .Q(\u2.mem[58][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13063_ (.D(_00942_),
    .CLK(clknet_leaf_48_clock),
    .Q(\u2.mem[58][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13064_ (.D(_00943_),
    .CLK(clknet_leaf_47_clock),
    .Q(\u2.mem[58][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13065_ (.D(_00944_),
    .CLK(clknet_leaf_47_clock),
    .Q(\u2.mem[58][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13066_ (.D(_00945_),
    .CLK(clknet_leaf_325_clock),
    .Q(\u2.mem[58][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13067_ (.D(_00946_),
    .CLK(clknet_leaf_248_clock),
    .Q(\u2.mem[59][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13068_ (.D(_00947_),
    .CLK(clknet_leaf_254_clock),
    .Q(\u2.mem[59][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13069_ (.D(_00948_),
    .CLK(clknet_leaf_259_clock),
    .Q(\u2.mem[59][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13070_ (.D(_00949_),
    .CLK(clknet_leaf_253_clock),
    .Q(\u2.mem[59][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13071_ (.D(_00950_),
    .CLK(clknet_leaf_240_clock),
    .Q(\u2.mem[59][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13072_ (.D(_00951_),
    .CLK(clknet_leaf_241_clock),
    .Q(\u2.mem[59][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13073_ (.D(_00952_),
    .CLK(clknet_leaf_236_clock),
    .Q(\u2.mem[59][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13074_ (.D(_00953_),
    .CLK(clknet_leaf_241_clock),
    .Q(\u2.mem[59][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13075_ (.D(_00954_),
    .CLK(clknet_leaf_25_clock),
    .Q(\u2.mem[59][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13076_ (.D(_00955_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u2.mem[59][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13077_ (.D(_00956_),
    .CLK(clknet_leaf_25_clock),
    .Q(\u2.mem[59][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13078_ (.D(_00957_),
    .CLK(clknet_leaf_25_clock),
    .Q(\u2.mem[59][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13079_ (.D(_00958_),
    .CLK(clknet_leaf_43_clock),
    .Q(\u2.mem[59][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13080_ (.D(_00959_),
    .CLK(clknet_leaf_43_clock),
    .Q(\u2.mem[59][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13081_ (.D(_00960_),
    .CLK(clknet_leaf_40_clock),
    .Q(\u2.mem[59][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13082_ (.D(_00961_),
    .CLK(clknet_leaf_42_clock),
    .Q(\u2.mem[59][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13083_ (.D(_00962_),
    .CLK(clknet_leaf_267_clock),
    .Q(\u2.mem[60][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13084_ (.D(_00963_),
    .CLK(clknet_leaf_261_clock),
    .Q(\u2.mem[60][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13085_ (.D(_00964_),
    .CLK(clknet_leaf_260_clock),
    .Q(\u2.mem[60][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13086_ (.D(_00965_),
    .CLK(clknet_leaf_267_clock),
    .Q(\u2.mem[60][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13087_ (.D(_00966_),
    .CLK(clknet_leaf_245_clock),
    .Q(\u2.mem[60][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13088_ (.D(_00967_),
    .CLK(clknet_leaf_245_clock),
    .Q(\u2.mem[60][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13089_ (.D(_00968_),
    .CLK(clknet_leaf_241_clock),
    .Q(\u2.mem[60][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13090_ (.D(_00969_),
    .CLK(clknet_leaf_242_clock),
    .Q(\u2.mem[60][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13091_ (.D(_00970_),
    .CLK(clknet_leaf_22_clock),
    .Q(\u2.mem[60][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13092_ (.D(_00971_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u2.mem[60][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13093_ (.D(_00972_),
    .CLK(clknet_leaf_24_clock),
    .Q(\u2.mem[60][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13094_ (.D(_00973_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u2.mem[60][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13095_ (.D(_00974_),
    .CLK(clknet_leaf_46_clock),
    .Q(\u2.mem[60][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13096_ (.D(_00975_),
    .CLK(clknet_leaf_47_clock),
    .Q(\u2.mem[60][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13097_ (.D(_00976_),
    .CLK(clknet_leaf_45_clock),
    .Q(\u2.mem[60][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13098_ (.D(_00977_),
    .CLK(clknet_leaf_45_clock),
    .Q(\u2.mem[60][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13099_ (.D(_00978_),
    .CLK(clknet_leaf_245_clock),
    .Q(\u2.mem[61][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13100_ (.D(_00979_),
    .CLK(clknet_leaf_264_clock),
    .Q(\u2.mem[61][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13101_ (.D(_00980_),
    .CLK(clknet_leaf_266_clock),
    .Q(\u2.mem[61][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13102_ (.D(_00981_),
    .CLK(clknet_leaf_266_clock),
    .Q(\u2.mem[61][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13103_ (.D(_00982_),
    .CLK(clknet_leaf_312_clock),
    .Q(\u2.mem[61][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13104_ (.D(_00983_),
    .CLK(clknet_leaf_243_clock),
    .Q(\u2.mem[61][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13105_ (.D(_00984_),
    .CLK(clknet_leaf_314_clock),
    .Q(\u2.mem[61][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13106_ (.D(_00985_),
    .CLK(clknet_leaf_241_clock),
    .Q(\u2.mem[61][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13107_ (.D(_00986_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u2.mem[61][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13108_ (.D(_00987_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u2.mem[61][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13109_ (.D(_00988_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u2.mem[61][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13110_ (.D(_00989_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u2.mem[61][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13111_ (.D(_00990_),
    .CLK(clknet_leaf_38_clock),
    .Q(\u2.mem[61][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13112_ (.D(_00991_),
    .CLK(clknet_leaf_39_clock),
    .Q(\u2.mem[61][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13113_ (.D(_00992_),
    .CLK(clknet_leaf_327_clock),
    .Q(\u2.mem[61][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13114_ (.D(_00993_),
    .CLK(clknet_leaf_333_clock),
    .Q(\u2.mem[61][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13115_ (.D(_00994_),
    .CLK(clknet_5_22_0_clock),
    .Q(\u2.mem[62][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13116_ (.D(_00995_),
    .CLK(clknet_leaf_261_clock),
    .Q(\u2.mem[62][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13117_ (.D(_00996_),
    .CLK(clknet_leaf_261_clock),
    .Q(\u2.mem[62][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13118_ (.D(_00997_),
    .CLK(clknet_leaf_266_clock),
    .Q(\u2.mem[62][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13119_ (.D(_00998_),
    .CLK(clknet_leaf_243_clock),
    .Q(\u2.mem[62][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13120_ (.D(_00999_),
    .CLK(clknet_leaf_244_clock),
    .Q(\u2.mem[62][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13121_ (.D(_01000_),
    .CLK(clknet_leaf_314_clock),
    .Q(\u2.mem[62][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13122_ (.D(_01001_),
    .CLK(clknet_leaf_242_clock),
    .Q(\u2.mem[62][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13123_ (.D(_01002_),
    .CLK(clknet_leaf_21_clock),
    .Q(\u2.mem[62][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13124_ (.D(_01003_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u2.mem[62][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13125_ (.D(_01004_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u2.mem[62][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13126_ (.D(_01005_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u2.mem[62][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13127_ (.D(_01006_),
    .CLK(clknet_leaf_327_clock),
    .Q(\u2.mem[62][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13128_ (.D(_01007_),
    .CLK(clknet_leaf_46_clock),
    .Q(\u2.mem[62][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13129_ (.D(_01008_),
    .CLK(clknet_leaf_327_clock),
    .Q(\u2.mem[62][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13130_ (.D(_01009_),
    .CLK(clknet_leaf_327_clock),
    .Q(\u2.mem[62][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13131_ (.D(_01010_),
    .CLK(clknet_leaf_246_clock),
    .Q(\u2.mem[63][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13132_ (.D(_01011_),
    .CLK(clknet_leaf_267_clock),
    .Q(\u2.mem[63][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13133_ (.D(_01012_),
    .CLK(clknet_leaf_268_clock),
    .Q(\u2.mem[63][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13134_ (.D(_01013_),
    .CLK(clknet_leaf_268_clock),
    .Q(\u2.mem[63][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13135_ (.D(_01014_),
    .CLK(clknet_leaf_314_clock),
    .Q(\u2.mem[63][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13136_ (.D(_01015_),
    .CLK(clknet_leaf_315_clock),
    .Q(\u2.mem[63][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13137_ (.D(_01016_),
    .CLK(clknet_leaf_315_clock),
    .Q(\u2.mem[63][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13138_ (.D(_01017_),
    .CLK(clknet_leaf_314_clock),
    .Q(\u2.mem[63][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13139_ (.D(_01018_),
    .CLK(clknet_leaf_21_clock),
    .Q(\u2.mem[63][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13140_ (.D(_01019_),
    .CLK(clknet_leaf_22_clock),
    .Q(\u2.mem[63][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13141_ (.D(_01020_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u2.mem[63][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13142_ (.D(_01021_),
    .CLK(clknet_leaf_23_clock),
    .Q(\u2.mem[63][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13143_ (.D(_01022_),
    .CLK(clknet_leaf_39_clock),
    .Q(\u2.mem[63][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13144_ (.D(_01023_),
    .CLK(clknet_leaf_39_clock),
    .Q(\u2.mem[63][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13145_ (.D(_01024_),
    .CLK(clknet_leaf_39_clock),
    .Q(\u2.mem[63][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13146_ (.D(_01025_),
    .CLK(clknet_leaf_38_clock),
    .Q(\u2.mem[63][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13147_ (.D(_01026_),
    .CLK(clknet_leaf_265_clock),
    .Q(\u2.mem[128][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13148_ (.D(_01027_),
    .CLK(clknet_leaf_263_clock),
    .Q(\u2.mem[128][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13149_ (.D(_01028_),
    .CLK(clknet_leaf_264_clock),
    .Q(\u2.mem[128][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13150_ (.D(_01029_),
    .CLK(clknet_leaf_262_clock),
    .Q(\u2.mem[128][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13151_ (.D(_01030_),
    .CLK(clknet_leaf_269_clock),
    .Q(\u2.mem[128][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13152_ (.D(_01031_),
    .CLK(clknet_leaf_245_clock),
    .Q(\u2.mem[128][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13153_ (.D(_01032_),
    .CLK(clknet_leaf_268_clock),
    .Q(\u2.mem[129][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13154_ (.D(_01033_),
    .CLK(clknet_leaf_263_clock),
    .Q(\u2.mem[129][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13155_ (.D(_01034_),
    .CLK(clknet_leaf_261_clock),
    .Q(\u2.mem[129][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13156_ (.D(_01035_),
    .CLK(clknet_leaf_262_clock),
    .Q(\u2.mem[129][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13157_ (.D(_01036_),
    .CLK(clknet_leaf_269_clock),
    .Q(\u2.mem[129][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13158_ (.D(_01037_),
    .CLK(clknet_leaf_269_clock),
    .Q(\u2.mem[129][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13159_ (.D(_01038_),
    .CLK(clknet_leaf_274_clock),
    .Q(\u2.mem[130][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13160_ (.D(_01039_),
    .CLK(clknet_leaf_276_clock),
    .Q(\u2.mem[130][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13161_ (.D(_01040_),
    .CLK(clknet_leaf_276_clock),
    .Q(\u2.mem[130][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13162_ (.D(_01041_),
    .CLK(clknet_leaf_275_clock),
    .Q(\u2.mem[130][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13163_ (.D(_01042_),
    .CLK(clknet_leaf_274_clock),
    .Q(\u2.mem[130][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13164_ (.D(_01043_),
    .CLK(clknet_leaf_270_clock),
    .Q(\u2.mem[130][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13165_ (.D(_01044_),
    .CLK(clknet_leaf_264_clock),
    .Q(\u2.mem[131][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13166_ (.D(_01045_),
    .CLK(clknet_leaf_263_clock),
    .Q(\u2.mem[131][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13167_ (.D(_01046_),
    .CLK(clknet_leaf_263_clock),
    .Q(\u2.mem[131][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13168_ (.D(_01047_),
    .CLK(clknet_leaf_263_clock),
    .Q(\u2.mem[131][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13169_ (.D(_01048_),
    .CLK(clknet_leaf_265_clock),
    .Q(\u2.mem[131][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13170_ (.D(_01049_),
    .CLK(clknet_leaf_268_clock),
    .Q(\u2.mem[131][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13171_ (.D(_01050_),
    .CLK(clknet_leaf_264_clock),
    .Q(\u2.mem[132][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13172_ (.D(_01051_),
    .CLK(clknet_leaf_263_clock),
    .Q(\u2.mem[132][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13173_ (.D(_01052_),
    .CLK(clknet_leaf_263_clock),
    .Q(\u2.mem[132][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13174_ (.D(_01053_),
    .CLK(clknet_leaf_275_clock),
    .Q(\u2.mem[132][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13175_ (.D(_01054_),
    .CLK(clknet_leaf_265_clock),
    .Q(\u2.mem[132][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13176_ (.D(_01055_),
    .CLK(clknet_leaf_269_clock),
    .Q(\u2.mem[132][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13177_ (.D(_01056_),
    .CLK(clknet_leaf_275_clock),
    .Q(\u2.mem[133][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13178_ (.D(_01057_),
    .CLK(clknet_leaf_276_clock),
    .Q(\u2.mem[133][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13179_ (.D(_01058_),
    .CLK(clknet_leaf_275_clock),
    .Q(\u2.mem[133][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13180_ (.D(_01059_),
    .CLK(clknet_leaf_275_clock),
    .Q(\u2.mem[133][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13181_ (.D(_01060_),
    .CLK(clknet_leaf_271_clock),
    .Q(\u2.mem[133][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13182_ (.D(_01061_),
    .CLK(clknet_leaf_271_clock),
    .Q(\u2.mem[133][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13183_ (.D(_01062_),
    .CLK(clknet_leaf_273_clock),
    .Q(\u2.mem[134][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13184_ (.D(_01063_),
    .CLK(clknet_leaf_277_clock),
    .Q(\u2.mem[134][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13185_ (.D(_01064_),
    .CLK(clknet_leaf_277_clock),
    .Q(\u2.mem[134][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13186_ (.D(_01065_),
    .CLK(clknet_leaf_276_clock),
    .Q(\u2.mem[134][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13187_ (.D(_01066_),
    .CLK(clknet_leaf_274_clock),
    .Q(\u2.mem[134][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13188_ (.D(_01067_),
    .CLK(clknet_leaf_270_clock),
    .Q(\u2.mem[134][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13189_ (.D(_01068_),
    .CLK(clknet_leaf_277_clock),
    .Q(\u2.mem[135][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13190_ (.D(_01069_),
    .CLK(clknet_leaf_279_clock),
    .Q(\u2.mem[135][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13191_ (.D(_01070_),
    .CLK(clknet_leaf_279_clock),
    .Q(\u2.mem[135][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13192_ (.D(_01071_),
    .CLK(clknet_leaf_276_clock),
    .Q(\u2.mem[135][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13193_ (.D(_01072_),
    .CLK(clknet_leaf_274_clock),
    .Q(\u2.mem[135][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13194_ (.D(_01073_),
    .CLK(clknet_leaf_272_clock),
    .Q(\u2.mem[135][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13195_ (.D(_01074_),
    .CLK(clknet_leaf_273_clock),
    .Q(\u2.mem[136][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13196_ (.D(_01075_),
    .CLK(clknet_leaf_277_clock),
    .Q(\u2.mem[136][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13197_ (.D(_01076_),
    .CLK(clknet_leaf_277_clock),
    .Q(\u2.mem[136][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13198_ (.D(_01077_),
    .CLK(clknet_leaf_276_clock),
    .Q(\u2.mem[136][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13199_ (.D(_01078_),
    .CLK(clknet_leaf_274_clock),
    .Q(\u2.mem[136][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13200_ (.D(_01079_),
    .CLK(clknet_leaf_271_clock),
    .Q(\u2.mem[136][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13201_ (.D(_01080_),
    .CLK(clknet_leaf_278_clock),
    .Q(\u2.mem[137][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13202_ (.D(_01081_),
    .CLK(clknet_leaf_280_clock),
    .Q(\u2.mem[137][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13203_ (.D(_01082_),
    .CLK(clknet_leaf_280_clock),
    .Q(\u2.mem[137][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13204_ (.D(_01083_),
    .CLK(clknet_leaf_276_clock),
    .Q(\u2.mem[137][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13205_ (.D(_01084_),
    .CLK(clknet_leaf_275_clock),
    .Q(\u2.mem[137][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13206_ (.D(_01085_),
    .CLK(clknet_leaf_271_clock),
    .Q(\u2.mem[137][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13207_ (.D(_01086_),
    .CLK(clknet_leaf_287_clock),
    .Q(\u2.mem[138][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13208_ (.D(_01087_),
    .CLK(clknet_leaf_281_clock),
    .Q(\u2.mem[138][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13209_ (.D(_01088_),
    .CLK(clknet_leaf_281_clock),
    .Q(\u2.mem[138][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13210_ (.D(_01089_),
    .CLK(clknet_leaf_281_clock),
    .Q(\u2.mem[138][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13211_ (.D(_01090_),
    .CLK(clknet_leaf_287_clock),
    .Q(\u2.mem[138][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13212_ (.D(_01091_),
    .CLK(clknet_leaf_291_clock),
    .Q(\u2.mem[138][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13213_ (.D(_01092_),
    .CLK(clknet_leaf_282_clock),
    .Q(\u2.mem[139][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13214_ (.D(_01093_),
    .CLK(clknet_leaf_282_clock),
    .Q(\u2.mem[139][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13215_ (.D(_01094_),
    .CLK(clknet_leaf_283_clock),
    .Q(\u2.mem[139][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13216_ (.D(_01095_),
    .CLK(clknet_leaf_282_clock),
    .Q(\u2.mem[139][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13217_ (.D(_01096_),
    .CLK(clknet_leaf_286_clock),
    .Q(\u2.mem[139][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13218_ (.D(_01097_),
    .CLK(clknet_leaf_283_clock),
    .Q(\u2.mem[139][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13219_ (.D(_01098_),
    .CLK(clknet_leaf_283_clock),
    .Q(\u2.mem[140][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13220_ (.D(_01099_),
    .CLK(clknet_leaf_282_clock),
    .Q(\u2.mem[140][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13221_ (.D(_01100_),
    .CLK(clknet_leaf_281_clock),
    .Q(\u2.mem[140][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13222_ (.D(_01101_),
    .CLK(clknet_leaf_280_clock),
    .Q(\u2.mem[140][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13223_ (.D(_01102_),
    .CLK(clknet_leaf_286_clock),
    .Q(\u2.mem[140][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13224_ (.D(_01103_),
    .CLK(clknet_leaf_286_clock),
    .Q(\u2.mem[140][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13225_ (.D(_01104_),
    .CLK(clknet_leaf_283_clock),
    .Q(\u2.mem[141][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13226_ (.D(_01105_),
    .CLK(clknet_leaf_279_clock),
    .Q(\u2.mem[141][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13227_ (.D(_01106_),
    .CLK(clknet_leaf_279_clock),
    .Q(\u2.mem[141][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13228_ (.D(_01107_),
    .CLK(clknet_leaf_280_clock),
    .Q(\u2.mem[141][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13229_ (.D(_01108_),
    .CLK(clknet_leaf_286_clock),
    .Q(\u2.mem[141][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13230_ (.D(_01109_),
    .CLK(clknet_leaf_279_clock),
    .Q(\u2.mem[141][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13231_ (.D(_01110_),
    .CLK(clknet_leaf_284_clock),
    .Q(\u2.mem[142][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13232_ (.D(_01111_),
    .CLK(clknet_leaf_279_clock),
    .Q(\u2.mem[142][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13233_ (.D(_01112_),
    .CLK(clknet_leaf_285_clock),
    .Q(\u2.mem[142][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13234_ (.D(_01113_),
    .CLK(clknet_leaf_278_clock),
    .Q(\u2.mem[142][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13235_ (.D(_01114_),
    .CLK(clknet_leaf_272_clock),
    .Q(\u2.mem[142][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13236_ (.D(_01115_),
    .CLK(clknet_leaf_273_clock),
    .Q(\u2.mem[142][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13237_ (.D(_01116_),
    .CLK(clknet_leaf_284_clock),
    .Q(\u2.mem[143][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13238_ (.D(_01117_),
    .CLK(clknet_leaf_284_clock),
    .Q(\u2.mem[143][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13239_ (.D(_01118_),
    .CLK(clknet_leaf_284_clock),
    .Q(\u2.mem[143][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13240_ (.D(_01119_),
    .CLK(clknet_leaf_278_clock),
    .Q(\u2.mem[143][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13241_ (.D(_01120_),
    .CLK(clknet_leaf_272_clock),
    .Q(\u2.mem[143][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13242_ (.D(_01121_),
    .CLK(clknet_leaf_278_clock),
    .Q(\u2.mem[143][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13243_ (.D(_01122_),
    .CLK(clknet_leaf_291_clock),
    .Q(\u2.mem[144][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13244_ (.D(_01123_),
    .CLK(clknet_leaf_291_clock),
    .Q(\u2.mem[144][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13245_ (.D(_01124_),
    .CLK(clknet_leaf_285_clock),
    .Q(\u2.mem[144][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13246_ (.D(_01125_),
    .CLK(clknet_leaf_272_clock),
    .Q(\u2.mem[144][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13247_ (.D(_01126_),
    .CLK(clknet_leaf_272_clock),
    .Q(\u2.mem[144][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13248_ (.D(_01127_),
    .CLK(clknet_leaf_272_clock),
    .Q(\u2.mem[144][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13249_ (.D(_01128_),
    .CLK(clknet_leaf_285_clock),
    .Q(\u2.mem[145][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13250_ (.D(_01129_),
    .CLK(clknet_leaf_285_clock),
    .Q(\u2.mem[145][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13251_ (.D(_01130_),
    .CLK(clknet_leaf_285_clock),
    .Q(\u2.mem[145][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13252_ (.D(_01131_),
    .CLK(clknet_leaf_291_clock),
    .Q(\u2.mem[145][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13253_ (.D(_01132_),
    .CLK(clknet_leaf_291_clock),
    .Q(\u2.mem[145][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13254_ (.D(_01133_),
    .CLK(clknet_leaf_291_clock),
    .Q(\u2.mem[145][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13255_ (.D(_01134_),
    .CLK(clknet_leaf_295_clock),
    .Q(\u2.mem[146][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13256_ (.D(_01135_),
    .CLK(clknet_leaf_311_clock),
    .Q(\u2.mem[146][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13257_ (.D(_01136_),
    .CLK(clknet_leaf_312_clock),
    .Q(\u2.mem[146][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13258_ (.D(_01137_),
    .CLK(clknet_leaf_312_clock),
    .Q(\u2.mem[146][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13259_ (.D(_01138_),
    .CLK(clknet_leaf_311_clock),
    .Q(\u2.mem[146][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13260_ (.D(_01139_),
    .CLK(clknet_leaf_295_clock),
    .Q(\u2.mem[146][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13261_ (.D(_01140_),
    .CLK(clknet_leaf_270_clock),
    .Q(\u2.mem[147][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13262_ (.D(_01141_),
    .CLK(clknet_leaf_271_clock),
    .Q(\u2.mem[147][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13263_ (.D(_01142_),
    .CLK(clknet_leaf_272_clock),
    .Q(\u2.mem[147][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13264_ (.D(_01143_),
    .CLK(clknet_leaf_270_clock),
    .Q(\u2.mem[147][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13265_ (.D(_01144_),
    .CLK(clknet_leaf_295_clock),
    .Q(\u2.mem[147][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13266_ (.D(_01145_),
    .CLK(clknet_leaf_295_clock),
    .Q(\u2.mem[147][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13267_ (.D(_01146_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u2.mem[148][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13268_ (.D(_01147_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u2.mem[148][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13269_ (.D(_01148_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u2.mem[148][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13270_ (.D(_01149_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u2.mem[148][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13271_ (.D(_01150_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u2.mem[148][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13272_ (.D(_01151_),
    .CLK(clknet_5_0_0_clock),
    .Q(\u2.mem[148][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13273_ (.D(_01152_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u2.mem[149][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13274_ (.D(_01153_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u2.mem[149][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13275_ (.D(_01154_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u2.mem[149][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13276_ (.D(_01155_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u2.mem[149][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13277_ (.D(_01156_),
    .CLK(clknet_leaf_10_clock),
    .Q(\u2.mem[149][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13278_ (.D(_01157_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u2.mem[149][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13279_ (.D(_01158_),
    .CLK(clknet_leaf_361_clock),
    .Q(\u2.mem[150][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13280_ (.D(_01159_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u2.mem[150][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13281_ (.D(_01160_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u2.mem[150][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13282_ (.D(_01161_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u2.mem[150][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13283_ (.D(_01162_),
    .CLK(clknet_leaf_360_clock),
    .Q(\u2.mem[150][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13284_ (.D(_01163_),
    .CLK(clknet_leaf_1_clock),
    .Q(\u2.mem[150][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13285_ (.D(_01164_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u2.mem[151][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13286_ (.D(_01165_),
    .CLK(clknet_leaf_1_clock),
    .Q(\u2.mem[151][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13287_ (.D(_01166_),
    .CLK(clknet_leaf_364_clock),
    .Q(\u2.mem[151][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13288_ (.D(_01167_),
    .CLK(clknet_leaf_364_clock),
    .Q(\u2.mem[151][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13289_ (.D(_01168_),
    .CLK(clknet_leaf_1_clock),
    .Q(\u2.mem[151][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13290_ (.D(_01169_),
    .CLK(clknet_leaf_354_clock),
    .Q(\u2.mem[151][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13291_ (.D(_01170_),
    .CLK(clknet_leaf_361_clock),
    .Q(\u2.mem[152][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13292_ (.D(_01171_),
    .CLK(clknet_leaf_0_clock),
    .Q(\u2.mem[152][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13293_ (.D(_01172_),
    .CLK(clknet_leaf_364_clock),
    .Q(\u2.mem[152][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13294_ (.D(_01173_),
    .CLK(clknet_leaf_364_clock),
    .Q(\u2.mem[152][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13295_ (.D(_01174_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u2.mem[152][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13296_ (.D(_01175_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u2.mem[152][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13297_ (.D(_01176_),
    .CLK(clknet_leaf_363_clock),
    .Q(\u2.mem[153][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13298_ (.D(_01177_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u2.mem[153][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13299_ (.D(_01178_),
    .CLK(clknet_leaf_363_clock),
    .Q(\u2.mem[153][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13300_ (.D(_01179_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u2.mem[153][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13301_ (.D(_01180_),
    .CLK(clknet_leaf_2_clock),
    .Q(\u2.mem[153][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13302_ (.D(_01181_),
    .CLK(clknet_leaf_7_clock),
    .Q(\u2.mem[153][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13303_ (.D(_01182_),
    .CLK(clknet_leaf_362_clock),
    .Q(\u2.mem[154][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13304_ (.D(_01183_),
    .CLK(clknet_leaf_362_clock),
    .Q(\u2.mem[154][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13305_ (.D(_01184_),
    .CLK(clknet_leaf_358_clock),
    .Q(\u2.mem[154][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13306_ (.D(_01185_),
    .CLK(clknet_leaf_358_clock),
    .Q(\u2.mem[154][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13307_ (.D(_01186_),
    .CLK(clknet_leaf_359_clock),
    .Q(\u2.mem[154][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13308_ (.D(_01187_),
    .CLK(clknet_leaf_353_clock),
    .Q(\u2.mem[154][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13309_ (.D(_01188_),
    .CLK(clknet_leaf_348_clock),
    .Q(\u2.mem[155][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13310_ (.D(_01189_),
    .CLK(clknet_leaf_348_clock),
    .Q(\u2.mem[155][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13311_ (.D(_01190_),
    .CLK(clknet_leaf_347_clock),
    .Q(\u2.mem[155][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13312_ (.D(_01191_),
    .CLK(clknet_leaf_348_clock),
    .Q(\u2.mem[155][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13313_ (.D(_01192_),
    .CLK(clknet_leaf_349_clock),
    .Q(\u2.mem[155][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13314_ (.D(_01193_),
    .CLK(clknet_leaf_349_clock),
    .Q(\u2.mem[155][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13315_ (.D(_01194_),
    .CLK(clknet_leaf_300_clock),
    .Q(\u2.mem[156][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13316_ (.D(_01195_),
    .CLK(clknet_leaf_300_clock),
    .Q(\u2.mem[156][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13317_ (.D(_01196_),
    .CLK(clknet_leaf_301_clock),
    .Q(\u2.mem[156][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13318_ (.D(_01197_),
    .CLK(clknet_leaf_301_clock),
    .Q(\u2.mem[156][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13319_ (.D(_01198_),
    .CLK(clknet_leaf_301_clock),
    .Q(\u2.mem[156][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13320_ (.D(_01199_),
    .CLK(clknet_leaf_306_clock),
    .Q(\u2.mem[156][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13321_ (.D(_01200_),
    .CLK(clknet_leaf_303_clock),
    .Q(\u2.mem[157][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13322_ (.D(_01201_),
    .CLK(clknet_leaf_342_clock),
    .Q(\u2.mem[157][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13323_ (.D(_01202_),
    .CLK(clknet_leaf_303_clock),
    .Q(\u2.mem[157][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13324_ (.D(_01203_),
    .CLK(clknet_leaf_342_clock),
    .Q(\u2.mem[157][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13325_ (.D(_01204_),
    .CLK(clknet_leaf_342_clock),
    .Q(\u2.mem[157][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13326_ (.D(_01205_),
    .CLK(clknet_leaf_304_clock),
    .Q(\u2.mem[157][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13327_ (.D(_01206_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u2.mem[158][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13328_ (.D(_01207_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u2.mem[158][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13329_ (.D(_01208_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u2.mem[158][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13330_ (.D(_01209_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u2.mem[158][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13331_ (.D(_01210_),
    .CLK(clknet_leaf_353_clock),
    .Q(\u2.mem[158][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13332_ (.D(_01211_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u2.mem[158][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13333_ (.D(_01212_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u2.mem[159][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13334_ (.D(_01213_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u2.mem[159][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13335_ (.D(_01214_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u2.mem[159][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13336_ (.D(_01215_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u2.mem[159][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13337_ (.D(_01216_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u2.mem[159][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13338_ (.D(_01217_),
    .CLK(clknet_leaf_9_clock),
    .Q(\u2.mem[159][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13339_ (.D(_01218_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u2.mem[160][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13340_ (.D(_01219_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u2.mem[160][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13341_ (.D(_01220_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u2.mem[160][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13342_ (.D(_01221_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u2.mem[160][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13343_ (.D(_01222_),
    .CLK(clknet_leaf_3_clock),
    .Q(\u2.mem[160][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13344_ (.D(_01223_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u2.mem[160][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13345_ (.D(_01224_),
    .CLK(clknet_leaf_4_clock),
    .Q(\u2.mem[161][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13346_ (.D(_01225_),
    .CLK(clknet_leaf_5_clock),
    .Q(\u2.mem[161][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13347_ (.D(_01226_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u2.mem[161][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13348_ (.D(_01227_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u2.mem[161][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13349_ (.D(_01228_),
    .CLK(clknet_leaf_10_clock),
    .Q(\u2.mem[161][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13350_ (.D(_01229_),
    .CLK(clknet_leaf_8_clock),
    .Q(\u2.mem[161][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13351_ (.D(_01230_),
    .CLK(clknet_leaf_361_clock),
    .Q(\u2.mem[162][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13352_ (.D(_01231_),
    .CLK(clknet_leaf_361_clock),
    .Q(\u2.mem[162][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13353_ (.D(_01232_),
    .CLK(clknet_leaf_358_clock),
    .Q(\u2.mem[162][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13354_ (.D(_01233_),
    .CLK(clknet_leaf_359_clock),
    .Q(\u2.mem[162][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13355_ (.D(_01234_),
    .CLK(clknet_leaf_360_clock),
    .Q(\u2.mem[162][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13356_ (.D(_01235_),
    .CLK(clknet_leaf_360_clock),
    .Q(\u2.mem[162][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13357_ (.D(_01236_),
    .CLK(clknet_leaf_356_clock),
    .Q(\u2.mem[163][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13358_ (.D(_01237_),
    .CLK(clknet_leaf_356_clock),
    .Q(\u2.mem[163][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13359_ (.D(_01238_),
    .CLK(clknet_leaf_357_clock),
    .Q(\u2.mem[163][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13360_ (.D(_01239_),
    .CLK(clknet_leaf_356_clock),
    .Q(\u2.mem[163][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13361_ (.D(_01240_),
    .CLK(clknet_leaf_355_clock),
    .Q(\u2.mem[163][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13362_ (.D(_01241_),
    .CLK(clknet_leaf_354_clock),
    .Q(\u2.mem[163][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13363_ (.D(_01242_),
    .CLK(clknet_leaf_358_clock),
    .Q(\u2.mem[164][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13364_ (.D(_01243_),
    .CLK(clknet_leaf_358_clock),
    .Q(\u2.mem[164][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13365_ (.D(_01244_),
    .CLK(clknet_leaf_358_clock),
    .Q(\u2.mem[164][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13366_ (.D(_01245_),
    .CLK(clknet_leaf_359_clock),
    .Q(\u2.mem[164][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13367_ (.D(_01246_),
    .CLK(clknet_leaf_354_clock),
    .Q(\u2.mem[164][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13368_ (.D(_01247_),
    .CLK(clknet_leaf_359_clock),
    .Q(\u2.mem[164][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13369_ (.D(_01248_),
    .CLK(clknet_leaf_356_clock),
    .Q(\u2.mem[165][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13370_ (.D(_01249_),
    .CLK(clknet_leaf_357_clock),
    .Q(\u2.mem[165][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13371_ (.D(_01250_),
    .CLK(clknet_leaf_357_clock),
    .Q(\u2.mem[165][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13372_ (.D(_01251_),
    .CLK(clknet_leaf_359_clock),
    .Q(\u2.mem[165][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13373_ (.D(_01252_),
    .CLK(clknet_leaf_354_clock),
    .Q(\u2.mem[165][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13374_ (.D(_01253_),
    .CLK(clknet_leaf_355_clock),
    .Q(\u2.mem[165][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13375_ (.D(_01254_),
    .CLK(clknet_leaf_352_clock),
    .Q(\u2.mem[166][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13376_ (.D(_01255_),
    .CLK(clknet_leaf_10_clock),
    .Q(\u2.mem[166][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13377_ (.D(_01256_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u2.mem[166][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13378_ (.D(_01257_),
    .CLK(clknet_leaf_36_clock),
    .Q(\u2.mem[166][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13379_ (.D(_01258_),
    .CLK(clknet_leaf_352_clock),
    .Q(\u2.mem[166][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13380_ (.D(_01259_),
    .CLK(clknet_leaf_352_clock),
    .Q(\u2.mem[166][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13381_ (.D(_01260_),
    .CLK(clknet_leaf_305_clock),
    .Q(\u2.mem[167][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13382_ (.D(_01261_),
    .CLK(clknet_leaf_309_clock),
    .Q(\u2.mem[167][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13383_ (.D(_01262_),
    .CLK(clknet_leaf_301_clock),
    .Q(\u2.mem[167][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13384_ (.D(_01263_),
    .CLK(clknet_leaf_301_clock),
    .Q(\u2.mem[167][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13385_ (.D(_01264_),
    .CLK(clknet_leaf_306_clock),
    .Q(\u2.mem[167][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13386_ (.D(_01265_),
    .CLK(clknet_leaf_306_clock),
    .Q(\u2.mem[167][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13387_ (.D(_01266_),
    .CLK(clknet_leaf_355_clock),
    .Q(\u2.mem[168][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13388_ (.D(_01267_),
    .CLK(clknet_leaf_355_clock),
    .Q(\u2.mem[168][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13389_ (.D(_01268_),
    .CLK(clknet_leaf_355_clock),
    .Q(\u2.mem[168][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13390_ (.D(_01269_),
    .CLK(clknet_leaf_355_clock),
    .Q(\u2.mem[168][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13391_ (.D(_01270_),
    .CLK(clknet_leaf_353_clock),
    .Q(\u2.mem[168][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13392_ (.D(_01271_),
    .CLK(clknet_leaf_353_clock),
    .Q(\u2.mem[168][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13393_ (.D(_01272_),
    .CLK(clknet_5_16_0_clock),
    .Q(\u2.mem[169][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13394_ (.D(_01273_),
    .CLK(clknet_leaf_310_clock),
    .Q(\u2.mem[169][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13395_ (.D(_01274_),
    .CLK(clknet_leaf_307_clock),
    .Q(\u2.mem[169][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13396_ (.D(_01275_),
    .CLK(clknet_leaf_310_clock),
    .Q(\u2.mem[169][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13397_ (.D(_01276_),
    .CLK(clknet_leaf_307_clock),
    .Q(\u2.mem[169][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13398_ (.D(_01277_),
    .CLK(clknet_leaf_307_clock),
    .Q(\u2.mem[169][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13399_ (.D(_01278_),
    .CLK(clknet_leaf_297_clock),
    .Q(\u2.mem[170][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13400_ (.D(_01279_),
    .CLK(clknet_leaf_301_clock),
    .Q(\u2.mem[170][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13401_ (.D(_01280_),
    .CLK(clknet_leaf_297_clock),
    .Q(\u2.mem[170][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13402_ (.D(_01281_),
    .CLK(clknet_leaf_298_clock),
    .Q(\u2.mem[170][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13403_ (.D(_01282_),
    .CLK(clknet_leaf_309_clock),
    .Q(\u2.mem[170][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13404_ (.D(_01283_),
    .CLK(clknet_leaf_305_clock),
    .Q(\u2.mem[170][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13405_ (.D(_01284_),
    .CLK(clknet_leaf_304_clock),
    .Q(\u2.mem[171][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13406_ (.D(_01285_),
    .CLK(clknet_leaf_304_clock),
    .Q(\u2.mem[171][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13407_ (.D(_01286_),
    .CLK(clknet_leaf_304_clock),
    .Q(\u2.mem[171][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13408_ (.D(_01287_),
    .CLK(clknet_leaf_304_clock),
    .Q(\u2.mem[171][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13409_ (.D(_01288_),
    .CLK(clknet_leaf_305_clock),
    .Q(\u2.mem[171][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13410_ (.D(_01289_),
    .CLK(clknet_leaf_305_clock),
    .Q(\u2.mem[171][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13411_ (.D(_01290_),
    .CLK(clknet_leaf_341_clock),
    .Q(\u2.mem[172][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13412_ (.D(_01291_),
    .CLK(clknet_leaf_344_clock),
    .Q(\u2.mem[172][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13413_ (.D(_01292_),
    .CLK(clknet_leaf_344_clock),
    .Q(\u2.mem[172][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13414_ (.D(_01293_),
    .CLK(clknet_leaf_342_clock),
    .Q(\u2.mem[172][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13415_ (.D(_01294_),
    .CLK(clknet_leaf_342_clock),
    .Q(\u2.mem[172][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13416_ (.D(_01295_),
    .CLK(clknet_leaf_341_clock),
    .Q(\u2.mem[172][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13417_ (.D(_01296_),
    .CLK(clknet_leaf_298_clock),
    .Q(\u2.mem[173][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13418_ (.D(_01297_),
    .CLK(clknet_leaf_299_clock),
    .Q(\u2.mem[173][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13419_ (.D(_01298_),
    .CLK(clknet_leaf_297_clock),
    .Q(\u2.mem[173][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13420_ (.D(_01299_),
    .CLK(clknet_leaf_298_clock),
    .Q(\u2.mem[173][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13421_ (.D(_01300_),
    .CLK(clknet_leaf_297_clock),
    .Q(\u2.mem[173][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13422_ (.D(_01301_),
    .CLK(clknet_leaf_309_clock),
    .Q(\u2.mem[173][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13423_ (.D(_01302_),
    .CLK(clknet_leaf_348_clock),
    .Q(\u2.mem[174][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13424_ (.D(_01303_),
    .CLK(clknet_leaf_347_clock),
    .Q(\u2.mem[174][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13425_ (.D(_01304_),
    .CLK(clknet_leaf_349_clock),
    .Q(\u2.mem[174][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13426_ (.D(_01305_),
    .CLK(clknet_leaf_349_clock),
    .Q(\u2.mem[174][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13427_ (.D(_01306_),
    .CLK(clknet_leaf_349_clock),
    .Q(\u2.mem[174][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13428_ (.D(_01307_),
    .CLK(clknet_leaf_350_clock),
    .Q(\u2.mem[174][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13429_ (.D(_01308_),
    .CLK(clknet_leaf_337_clock),
    .Q(\u2.mem[175][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13430_ (.D(_01309_),
    .CLK(clknet_5_4_0_clock),
    .Q(\u2.mem[175][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13431_ (.D(_01310_),
    .CLK(clknet_leaf_36_clock),
    .Q(\u2.mem[175][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13432_ (.D(_01311_),
    .CLK(clknet_leaf_336_clock),
    .Q(\u2.mem[175][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13433_ (.D(_01312_),
    .CLK(clknet_leaf_338_clock),
    .Q(\u2.mem[175][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13434_ (.D(_01313_),
    .CLK(clknet_leaf_337_clock),
    .Q(\u2.mem[175][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13435_ (.D(_01314_),
    .CLK(clknet_leaf_350_clock),
    .Q(\u2.mem[176][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13436_ (.D(_01315_),
    .CLK(clknet_leaf_350_clock),
    .Q(\u2.mem[176][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13437_ (.D(_01316_),
    .CLK(clknet_leaf_350_clock),
    .Q(\u2.mem[176][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13438_ (.D(_01317_),
    .CLK(clknet_5_5_0_clock),
    .Q(\u2.mem[176][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13439_ (.D(_01318_),
    .CLK(clknet_leaf_341_clock),
    .Q(\u2.mem[176][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13440_ (.D(_01319_),
    .CLK(clknet_leaf_341_clock),
    .Q(\u2.mem[176][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13441_ (.D(_01320_),
    .CLK(clknet_leaf_348_clock),
    .Q(\u2.mem[177][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13442_ (.D(_01321_),
    .CLK(clknet_leaf_356_clock),
    .Q(\u2.mem[177][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13443_ (.D(_01322_),
    .CLK(clknet_leaf_356_clock),
    .Q(\u2.mem[177][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13444_ (.D(_01323_),
    .CLK(clknet_leaf_349_clock),
    .Q(\u2.mem[177][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13445_ (.D(_01324_),
    .CLK(clknet_leaf_350_clock),
    .Q(\u2.mem[177][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13446_ (.D(_01325_),
    .CLK(clknet_leaf_350_clock),
    .Q(\u2.mem[177][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13447_ (.D(_01326_),
    .CLK(clknet_leaf_343_clock),
    .Q(\u2.mem[178][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13448_ (.D(_01327_),
    .CLK(clknet_leaf_343_clock),
    .Q(\u2.mem[178][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13449_ (.D(_01328_),
    .CLK(clknet_leaf_343_clock),
    .Q(\u2.mem[178][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13450_ (.D(_01329_),
    .CLK(clknet_leaf_343_clock),
    .Q(\u2.mem[178][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13451_ (.D(_01330_),
    .CLK(clknet_leaf_342_clock),
    .Q(\u2.mem[178][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13452_ (.D(_01331_),
    .CLK(clknet_leaf_342_clock),
    .Q(\u2.mem[178][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13453_ (.D(_01332_),
    .CLK(clknet_leaf_301_clock),
    .Q(\u2.mem[179][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13454_ (.D(_01333_),
    .CLK(clknet_leaf_300_clock),
    .Q(\u2.mem[179][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13455_ (.D(_01334_),
    .CLK(clknet_leaf_302_clock),
    .Q(\u2.mem[179][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13456_ (.D(_01335_),
    .CLK(clknet_leaf_304_clock),
    .Q(\u2.mem[179][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13457_ (.D(_01336_),
    .CLK(clknet_leaf_304_clock),
    .Q(\u2.mem[179][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13458_ (.D(_01337_),
    .CLK(clknet_leaf_306_clock),
    .Q(\u2.mem[179][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13459_ (.D(_01338_),
    .CLK(clknet_leaf_345_clock),
    .Q(\u2.mem[180][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13460_ (.D(_01339_),
    .CLK(clknet_leaf_345_clock),
    .Q(\u2.mem[180][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13461_ (.D(_01340_),
    .CLK(clknet_leaf_344_clock),
    .Q(\u2.mem[180][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13462_ (.D(_01341_),
    .CLK(clknet_leaf_346_clock),
    .Q(\u2.mem[180][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13463_ (.D(_01342_),
    .CLK(clknet_leaf_344_clock),
    .Q(\u2.mem[180][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13464_ (.D(_01343_),
    .CLK(clknet_leaf_344_clock),
    .Q(\u2.mem[180][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13465_ (.D(_01344_),
    .CLK(clknet_leaf_346_clock),
    .Q(\u2.mem[181][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13466_ (.D(_01345_),
    .CLK(clknet_leaf_347_clock),
    .Q(\u2.mem[181][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13467_ (.D(_01346_),
    .CLK(clknet_leaf_346_clock),
    .Q(\u2.mem[181][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13468_ (.D(_01347_),
    .CLK(clknet_leaf_346_clock),
    .Q(\u2.mem[181][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13469_ (.D(_01348_),
    .CLK(clknet_leaf_345_clock),
    .Q(\u2.mem[181][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13470_ (.D(_01349_),
    .CLK(clknet_leaf_347_clock),
    .Q(\u2.mem[181][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13471_ (.D(_01350_),
    .CLK(clknet_leaf_293_clock),
    .Q(\u2.mem[182][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13472_ (.D(_01351_),
    .CLK(clknet_leaf_294_clock),
    .Q(\u2.mem[182][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13473_ (.D(_01352_),
    .CLK(clknet_leaf_292_clock),
    .Q(\u2.mem[182][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13474_ (.D(_01353_),
    .CLK(clknet_leaf_293_clock),
    .Q(\u2.mem[182][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13475_ (.D(_01354_),
    .CLK(clknet_leaf_295_clock),
    .Q(\u2.mem[182][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13476_ (.D(_01355_),
    .CLK(clknet_leaf_295_clock),
    .Q(\u2.mem[182][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13477_ (.D(_01356_),
    .CLK(clknet_leaf_298_clock),
    .Q(\u2.mem[183][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13478_ (.D(_01357_),
    .CLK(clknet_leaf_290_clock),
    .Q(\u2.mem[183][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13479_ (.D(_01358_),
    .CLK(clknet_leaf_290_clock),
    .Q(\u2.mem[183][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13480_ (.D(_01359_),
    .CLK(clknet_leaf_289_clock),
    .Q(\u2.mem[183][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13481_ (.D(_01360_),
    .CLK(clknet_leaf_296_clock),
    .Q(\u2.mem[183][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13482_ (.D(_01361_),
    .CLK(clknet_leaf_298_clock),
    .Q(\u2.mem[183][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13483_ (.D(_01362_),
    .CLK(clknet_leaf_290_clock),
    .Q(\u2.mem[184][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13484_ (.D(_01363_),
    .CLK(clknet_leaf_290_clock),
    .Q(\u2.mem[184][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13485_ (.D(_01364_),
    .CLK(clknet_leaf_289_clock),
    .Q(\u2.mem[184][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13486_ (.D(_01365_),
    .CLK(clknet_leaf_298_clock),
    .Q(\u2.mem[184][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13487_ (.D(_01366_),
    .CLK(clknet_leaf_296_clock),
    .Q(\u2.mem[184][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13488_ (.D(_01367_),
    .CLK(clknet_leaf_298_clock),
    .Q(\u2.mem[184][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13489_ (.D(_01368_),
    .CLK(clknet_leaf_293_clock),
    .Q(\u2.mem[185][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13490_ (.D(_01369_),
    .CLK(clknet_leaf_292_clock),
    .Q(\u2.mem[185][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13491_ (.D(_01370_),
    .CLK(clknet_leaf_292_clock),
    .Q(\u2.mem[185][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13492_ (.D(_01371_),
    .CLK(clknet_leaf_292_clock),
    .Q(\u2.mem[185][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13493_ (.D(_01372_),
    .CLK(clknet_leaf_296_clock),
    .Q(\u2.mem[185][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13494_ (.D(_01373_),
    .CLK(clknet_leaf_295_clock),
    .Q(\u2.mem[185][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13495_ (.D(_01374_),
    .CLK(clknet_leaf_313_clock),
    .Q(\u2.mem[186][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13496_ (.D(_01375_),
    .CLK(clknet_leaf_312_clock),
    .Q(\u2.mem[186][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13497_ (.D(_01376_),
    .CLK(clknet_leaf_316_clock),
    .Q(\u2.mem[186][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13498_ (.D(_01377_),
    .CLK(clknet_leaf_313_clock),
    .Q(\u2.mem[186][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13499_ (.D(_01378_),
    .CLK(clknet_leaf_316_clock),
    .Q(\u2.mem[186][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13500_ (.D(_01379_),
    .CLK(clknet_leaf_317_clock),
    .Q(\u2.mem[186][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13501_ (.D(_01380_),
    .CLK(clknet_leaf_330_clock),
    .Q(\u2.mem[187][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13502_ (.D(_01381_),
    .CLK(clknet_leaf_331_clock),
    .Q(\u2.mem[187][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13503_ (.D(_01382_),
    .CLK(clknet_leaf_331_clock),
    .Q(\u2.mem[187][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13504_ (.D(_01383_),
    .CLK(clknet_leaf_331_clock),
    .Q(\u2.mem[187][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13505_ (.D(_01384_),
    .CLK(clknet_leaf_318_clock),
    .Q(\u2.mem[187][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13506_ (.D(_01385_),
    .CLK(clknet_leaf_330_clock),
    .Q(\u2.mem[187][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13507_ (.D(_01386_),
    .CLK(clknet_leaf_330_clock),
    .Q(\u2.mem[188][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13508_ (.D(_01387_),
    .CLK(clknet_leaf_331_clock),
    .Q(\u2.mem[188][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13509_ (.D(_01388_),
    .CLK(clknet_leaf_335_clock),
    .Q(\u2.mem[188][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13510_ (.D(_01389_),
    .CLK(clknet_leaf_335_clock),
    .Q(\u2.mem[188][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13511_ (.D(_01390_),
    .CLK(clknet_leaf_317_clock),
    .Q(\u2.mem[188][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13512_ (.D(_01391_),
    .CLK(clknet_leaf_330_clock),
    .Q(\u2.mem[188][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13513_ (.D(_01392_),
    .CLK(clknet_leaf_340_clock),
    .Q(\u2.mem[189][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13514_ (.D(_01393_),
    .CLK(clknet_leaf_340_clock),
    .Q(\u2.mem[189][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13515_ (.D(_01394_),
    .CLK(clknet_leaf_340_clock),
    .Q(\u2.mem[189][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13516_ (.D(_01395_),
    .CLK(clknet_leaf_338_clock),
    .Q(\u2.mem[189][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13517_ (.D(_01396_),
    .CLK(clknet_leaf_318_clock),
    .Q(\u2.mem[189][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13518_ (.D(_01397_),
    .CLK(clknet_leaf_330_clock),
    .Q(\u2.mem[189][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13519_ (.D(_01398_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u2.mem[190][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13520_ (.D(_01399_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u2.mem[190][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13521_ (.D(_01400_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u2.mem[190][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13522_ (.D(_01401_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u2.mem[190][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13523_ (.D(_01402_),
    .CLK(clknet_leaf_15_clock),
    .Q(\u2.mem[190][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13524_ (.D(_01403_),
    .CLK(clknet_leaf_15_clock),
    .Q(\u2.mem[190][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13525_ (.D(_01404_),
    .CLK(clknet_leaf_315_clock),
    .Q(\u2.mem[191][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13526_ (.D(_01405_),
    .CLK(clknet_leaf_314_clock),
    .Q(\u2.mem[191][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13527_ (.D(_01406_),
    .CLK(clknet_leaf_316_clock),
    .Q(\u2.mem[191][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13528_ (.D(_01407_),
    .CLK(clknet_leaf_317_clock),
    .Q(\u2.mem[191][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13529_ (.D(_01408_),
    .CLK(clknet_leaf_316_clock),
    .Q(\u2.mem[191][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13530_ (.D(_01409_),
    .CLK(clknet_leaf_317_clock),
    .Q(\u2.mem[191][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13531_ (.D(_01410_),
    .CLK(clknet_leaf_333_clock),
    .Q(\u2.mem[192][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13532_ (.D(_01411_),
    .CLK(clknet_leaf_334_clock),
    .Q(\u2.mem[192][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13533_ (.D(_01412_),
    .CLK(clknet_leaf_318_clock),
    .Q(\u2.mem[192][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13534_ (.D(_01413_),
    .CLK(clknet_leaf_318_clock),
    .Q(\u2.mem[192][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13535_ (.D(_01414_),
    .CLK(clknet_leaf_329_clock),
    .Q(\u2.mem[192][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13536_ (.D(_01415_),
    .CLK(clknet_leaf_318_clock),
    .Q(\u2.mem[192][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13537_ (.D(_01416_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u2.mem[192][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13538_ (.D(_01417_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u2.mem[192][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13539_ (.D(_01418_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u2.mem[192][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13540_ (.D(_01419_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u2.mem[192][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13541_ (.D(_01420_),
    .CLK(clknet_leaf_21_clock),
    .Q(\u2.mem[192][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13542_ (.D(_01421_),
    .CLK(clknet_leaf_21_clock),
    .Q(\u2.mem[192][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13543_ (.D(_01422_),
    .CLK(clknet_leaf_32_clock),
    .Q(\u2.mem[192][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13544_ (.D(_01423_),
    .CLK(clknet_leaf_32_clock),
    .Q(\u2.mem[192][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13545_ (.D(_01424_),
    .CLK(clknet_leaf_41_clock),
    .Q(\u2.mem[192][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13546_ (.D(_01425_),
    .CLK(clknet_leaf_38_clock),
    .Q(\u2.mem[192][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13547_ (.D(_01426_),
    .CLK(clknet_leaf_35_clock),
    .Q(\u2.mem[193][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13548_ (.D(_01427_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u2.mem[193][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13549_ (.D(_01428_),
    .CLK(clknet_leaf_11_clock),
    .Q(\u2.mem[193][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13550_ (.D(_01429_),
    .CLK(clknet_leaf_12_clock),
    .Q(\u2.mem[193][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13551_ (.D(_01430_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u2.mem[193][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13552_ (.D(_01431_),
    .CLK(clknet_leaf_13_clock),
    .Q(\u2.mem[193][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13553_ (.D(_01432_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u2.mem[193][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13554_ (.D(_01433_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u2.mem[193][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13555_ (.D(_01434_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u2.mem[193][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13556_ (.D(_01435_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u2.mem[193][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13557_ (.D(_01436_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u2.mem[193][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13558_ (.D(_01437_),
    .CLK(clknet_leaf_19_clock),
    .Q(\u2.mem[193][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13559_ (.D(_01438_),
    .CLK(clknet_leaf_33_clock),
    .Q(\u2.mem[193][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13560_ (.D(_01439_),
    .CLK(clknet_leaf_32_clock),
    .Q(\u2.mem[193][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13561_ (.D(_01440_),
    .CLK(clknet_leaf_32_clock),
    .Q(\u2.mem[193][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13562_ (.D(_01441_),
    .CLK(clknet_leaf_40_clock),
    .Q(\u2.mem[193][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13563_ (.D(_01442_),
    .CLK(clknet_leaf_16_clock),
    .Q(\u2.mem[194][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13564_ (.D(_01443_),
    .CLK(clknet_leaf_18_clock),
    .Q(\u2.mem[194][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13565_ (.D(_01444_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u2.mem[194][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13566_ (.D(_01445_),
    .CLK(clknet_leaf_17_clock),
    .Q(\u2.mem[194][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13567_ (.D(_01446_),
    .CLK(clknet_leaf_15_clock),
    .Q(\u2.mem[194][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13568_ (.D(_01447_),
    .CLK(clknet_leaf_15_clock),
    .Q(\u2.mem[194][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13569_ (.D(_01448_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u2.mem[194][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13570_ (.D(_01449_),
    .CLK(clknet_leaf_14_clock),
    .Q(\u2.mem[194][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13571_ (.D(_01450_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u2.mem[194][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13572_ (.D(_01451_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u2.mem[194][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13573_ (.D(_01452_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u2.mem[194][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13574_ (.D(_01453_),
    .CLK(clknet_leaf_20_clock),
    .Q(\u2.mem[194][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13575_ (.D(_01454_),
    .CLK(clknet_leaf_34_clock),
    .Q(\u2.mem[194][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13576_ (.D(_01455_),
    .CLK(clknet_leaf_32_clock),
    .Q(\u2.mem[194][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13577_ (.D(_01456_),
    .CLK(clknet_leaf_35_clock),
    .Q(\u2.mem[194][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13578_ (.D(_01457_),
    .CLK(clknet_leaf_37_clock),
    .Q(\u2.mem[194][15] ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(col_select_a[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(col_select_a[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(col_select_a[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(col_select_a[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(col_select_a[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(col_select_a[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(data_in_a[0]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(data_in_a[10]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(data_in_a[11]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(data_in_a[12]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(data_in_a[13]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(data_in_a[14]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(data_in_a[15]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(data_in_a[1]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(data_in_a[2]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(data_in_a[3]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(data_in_a[4]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(data_in_a[5]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(data_in_a[6]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(data_in_a[7]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(data_in_a[8]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(data_in_a[9]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(inverter_select_a),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(mem_address_a[0]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(mem_address_a[1]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(mem_address_a[2]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(mem_address_a[3]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(mem_address_a[4]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(mem_address_a[5]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(mem_address_a[6]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(mem_address_a[7]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(mem_address_a[8]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(mem_address_a[9]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(mem_write_n_a),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(output_active_a),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(row_col_select_a),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(row_select_a[0]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(row_select_a[1]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(row_select_a[2]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(row_select_a[3]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(row_select_a[4]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(row_select_a[5]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output43 (.I(net43),
    .Z(driver_io[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output44 (.I(net44),
    .Z(driver_io[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_clock (.I(clknet_5_0_0_clock),
    .Z(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_clock (.I(clknet_5_0_0_clock),
    .Z(clknet_leaf_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_clock (.I(clknet_5_0_0_clock),
    .Z(clknet_leaf_2_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_clock (.I(clknet_5_0_0_clock),
    .Z(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_clock (.I(clknet_5_0_0_clock),
    .Z(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_clock (.I(clknet_5_0_0_clock),
    .Z(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_clock (.I(clknet_5_0_0_clock),
    .Z(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_clock (.I(clknet_5_1_0_clock),
    .Z(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_clock (.I(clknet_5_1_0_clock),
    .Z(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_clock (.I(clknet_5_1_0_clock),
    .Z(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_clock (.I(clknet_5_3_0_clock),
    .Z(clknet_leaf_11_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_clock (.I(clknet_5_3_0_clock),
    .Z(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_clock (.I(clknet_5_3_0_clock),
    .Z(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_clock (.I(clknet_5_3_0_clock),
    .Z(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_clock (.I(clknet_5_2_0_clock),
    .Z(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_clock (.I(clknet_5_2_0_clock),
    .Z(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_clock (.I(clknet_5_2_0_clock),
    .Z(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_clock (.I(clknet_5_2_0_clock),
    .Z(clknet_leaf_18_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_clock (.I(clknet_5_2_0_clock),
    .Z(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_clock (.I(clknet_5_2_0_clock),
    .Z(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_clock (.I(clknet_5_2_0_clock),
    .Z(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_clock (.I(clknet_5_2_0_clock),
    .Z(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_clock (.I(clknet_5_2_0_clock),
    .Z(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_clock (.I(clknet_5_2_0_clock),
    .Z(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_clock (.I(clknet_5_2_0_clock),
    .Z(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_clock (.I(clknet_5_2_0_clock),
    .Z(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_clock (.I(clknet_5_2_0_clock),
    .Z(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_clock (.I(clknet_5_3_0_clock),
    .Z(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_clock (.I(clknet_5_3_0_clock),
    .Z(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_clock (.I(clknet_5_3_0_clock),
    .Z(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_clock (.I(clknet_5_3_0_clock),
    .Z(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_clock (.I(clknet_5_3_0_clock),
    .Z(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_clock (.I(clknet_5_3_0_clock),
    .Z(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_clock (.I(clknet_5_3_0_clock),
    .Z(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_clock (.I(clknet_5_3_0_clock),
    .Z(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_clock (.I(clknet_5_4_0_clock),
    .Z(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_clock (.I(clknet_5_6_0_clock),
    .Z(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_clock (.I(clknet_5_6_0_clock),
    .Z(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_clock (.I(clknet_5_6_0_clock),
    .Z(clknet_leaf_39_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_clock (.I(clknet_5_6_0_clock),
    .Z(clknet_leaf_40_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_clock (.I(clknet_5_6_0_clock),
    .Z(clknet_leaf_41_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_clock (.I(clknet_5_6_0_clock),
    .Z(clknet_leaf_42_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_clock (.I(clknet_5_6_0_clock),
    .Z(clknet_leaf_43_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_clock (.I(clknet_5_6_0_clock),
    .Z(clknet_leaf_44_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_clock (.I(clknet_5_6_0_clock),
    .Z(clknet_leaf_45_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_clock (.I(clknet_5_7_0_clock),
    .Z(clknet_leaf_46_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_clock (.I(clknet_5_7_0_clock),
    .Z(clknet_leaf_47_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_clock (.I(clknet_5_7_0_clock),
    .Z(clknet_leaf_48_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_clock (.I(clknet_5_7_0_clock),
    .Z(clknet_leaf_49_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_clock (.I(clknet_5_13_0_clock),
    .Z(clknet_leaf_50_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_clock (.I(clknet_5_13_0_clock),
    .Z(clknet_leaf_51_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_clock (.I(clknet_5_12_0_clock),
    .Z(clknet_leaf_52_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_clock (.I(clknet_5_12_0_clock),
    .Z(clknet_leaf_53_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_clock (.I(clknet_5_12_0_clock),
    .Z(clknet_leaf_54_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_clock (.I(clknet_5_12_0_clock),
    .Z(clknet_leaf_55_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_clock (.I(clknet_5_12_0_clock),
    .Z(clknet_leaf_56_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_clock (.I(clknet_5_12_0_clock),
    .Z(clknet_leaf_57_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_clock (.I(clknet_5_12_0_clock),
    .Z(clknet_leaf_58_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_clock (.I(clknet_5_12_0_clock),
    .Z(clknet_leaf_59_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_clock (.I(clknet_5_12_0_clock),
    .Z(clknet_leaf_60_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_clock (.I(clknet_5_9_0_clock),
    .Z(clknet_leaf_61_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_clock (.I(clknet_5_9_0_clock),
    .Z(clknet_leaf_62_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_clock (.I(clknet_5_9_0_clock),
    .Z(clknet_leaf_63_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_clock (.I(clknet_5_9_0_clock),
    .Z(clknet_leaf_64_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_clock (.I(clknet_5_9_0_clock),
    .Z(clknet_leaf_65_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_clock (.I(clknet_5_3_0_clock),
    .Z(clknet_leaf_66_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_clock (.I(clknet_5_9_0_clock),
    .Z(clknet_leaf_67_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_clock (.I(clknet_5_9_0_clock),
    .Z(clknet_leaf_68_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_clock (.I(clknet_5_9_0_clock),
    .Z(clknet_leaf_69_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_clock (.I(clknet_5_8_0_clock),
    .Z(clknet_leaf_70_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_clock (.I(clknet_5_8_0_clock),
    .Z(clknet_leaf_71_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_clock (.I(clknet_5_8_0_clock),
    .Z(clknet_leaf_72_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_clock (.I(clknet_5_8_0_clock),
    .Z(clknet_leaf_73_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_clock (.I(clknet_5_8_0_clock),
    .Z(clknet_leaf_74_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_clock (.I(clknet_5_8_0_clock),
    .Z(clknet_leaf_75_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_clock (.I(clknet_5_8_0_clock),
    .Z(clknet_leaf_76_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_clock (.I(clknet_5_8_0_clock),
    .Z(clknet_leaf_77_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_clock (.I(clknet_5_8_0_clock),
    .Z(clknet_leaf_78_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_clock (.I(clknet_5_8_0_clock),
    .Z(clknet_leaf_79_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_clock (.I(clknet_5_8_0_clock),
    .Z(clknet_leaf_80_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_clock (.I(clknet_5_8_0_clock),
    .Z(clknet_leaf_81_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_clock (.I(clknet_5_9_0_clock),
    .Z(clknet_leaf_82_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_clock (.I(clknet_5_9_0_clock),
    .Z(clknet_leaf_83_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_clock (.I(clknet_5_11_0_clock),
    .Z(clknet_leaf_84_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_clock (.I(clknet_5_11_0_clock),
    .Z(clknet_leaf_85_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_clock (.I(clknet_5_11_0_clock),
    .Z(clknet_leaf_86_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_clock (.I(clknet_5_11_0_clock),
    .Z(clknet_leaf_87_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_clock (.I(clknet_5_10_0_clock),
    .Z(clknet_leaf_88_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_clock (.I(clknet_5_10_0_clock),
    .Z(clknet_leaf_89_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_clock (.I(clknet_5_8_0_clock),
    .Z(clknet_leaf_90_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_clock (.I(clknet_5_10_0_clock),
    .Z(clknet_leaf_91_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_clock (.I(clknet_5_10_0_clock),
    .Z(clknet_leaf_92_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_clock (.I(clknet_5_10_0_clock),
    .Z(clknet_leaf_93_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_clock (.I(clknet_5_10_0_clock),
    .Z(clknet_leaf_94_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_clock (.I(clknet_5_10_0_clock),
    .Z(clknet_leaf_95_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_clock (.I(clknet_5_10_0_clock),
    .Z(clknet_leaf_96_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_clock (.I(clknet_5_10_0_clock),
    .Z(clknet_leaf_97_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_clock (.I(clknet_5_10_0_clock),
    .Z(clknet_leaf_98_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_clock (.I(clknet_5_10_0_clock),
    .Z(clknet_leaf_99_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_clock (.I(clknet_5_11_0_clock),
    .Z(clknet_leaf_100_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_clock (.I(clknet_5_11_0_clock),
    .Z(clknet_leaf_101_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_clock (.I(clknet_5_11_0_clock),
    .Z(clknet_leaf_102_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_clock (.I(clknet_5_11_0_clock),
    .Z(clknet_leaf_103_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_clock (.I(clknet_5_11_0_clock),
    .Z(clknet_leaf_104_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_clock (.I(clknet_5_11_0_clock),
    .Z(clknet_leaf_105_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_clock (.I(clknet_5_11_0_clock),
    .Z(clknet_leaf_106_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_clock (.I(clknet_5_11_0_clock),
    .Z(clknet_leaf_107_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_clock (.I(clknet_5_11_0_clock),
    .Z(clknet_leaf_108_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_clock (.I(clknet_5_11_0_clock),
    .Z(clknet_leaf_109_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_clock (.I(clknet_5_14_0_clock),
    .Z(clknet_leaf_110_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_111_clock (.I(clknet_5_14_0_clock),
    .Z(clknet_leaf_111_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_clock (.I(clknet_5_14_0_clock),
    .Z(clknet_leaf_112_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_113_clock (.I(clknet_5_14_0_clock),
    .Z(clknet_leaf_113_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_clock (.I(clknet_5_14_0_clock),
    .Z(clknet_leaf_114_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_clock (.I(clknet_5_14_0_clock),
    .Z(clknet_leaf_115_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_116_clock (.I(clknet_5_14_0_clock),
    .Z(clknet_leaf_116_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_clock (.I(clknet_5_14_0_clock),
    .Z(clknet_leaf_117_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_118_clock (.I(clknet_5_15_0_clock),
    .Z(clknet_leaf_118_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_119_clock (.I(clknet_5_15_0_clock),
    .Z(clknet_leaf_119_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_120_clock (.I(clknet_5_15_0_clock),
    .Z(clknet_leaf_120_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_121_clock (.I(clknet_5_15_0_clock),
    .Z(clknet_leaf_121_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_122_clock (.I(clknet_5_15_0_clock),
    .Z(clknet_leaf_122_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_123_clock (.I(clknet_5_15_0_clock),
    .Z(clknet_leaf_123_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_124_clock (.I(clknet_5_15_0_clock),
    .Z(clknet_leaf_124_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_125_clock (.I(clknet_5_15_0_clock),
    .Z(clknet_leaf_125_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_126_clock (.I(clknet_5_15_0_clock),
    .Z(clknet_leaf_126_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_127_clock (.I(clknet_5_15_0_clock),
    .Z(clknet_leaf_127_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_128_clock (.I(clknet_5_14_0_clock),
    .Z(clknet_leaf_128_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_129_clock (.I(clknet_5_14_0_clock),
    .Z(clknet_leaf_129_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_130_clock (.I(clknet_5_14_0_clock),
    .Z(clknet_leaf_130_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_131_clock (.I(clknet_5_12_0_clock),
    .Z(clknet_leaf_131_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_132_clock (.I(clknet_5_12_0_clock),
    .Z(clknet_leaf_132_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_133_clock (.I(clknet_5_12_0_clock),
    .Z(clknet_leaf_133_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_134_clock (.I(clknet_5_12_0_clock),
    .Z(clknet_leaf_134_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_135_clock (.I(clknet_5_13_0_clock),
    .Z(clknet_leaf_135_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_136_clock (.I(clknet_5_13_0_clock),
    .Z(clknet_leaf_136_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_137_clock (.I(clknet_5_13_0_clock),
    .Z(clknet_leaf_137_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_138_clock (.I(clknet_5_13_0_clock),
    .Z(clknet_leaf_138_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_139_clock (.I(clknet_5_13_0_clock),
    .Z(clknet_leaf_139_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_140_clock (.I(clknet_5_13_0_clock),
    .Z(clknet_leaf_140_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_141_clock (.I(clknet_5_13_0_clock),
    .Z(clknet_leaf_141_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_143_clock (.I(clknet_5_24_0_clock),
    .Z(clknet_leaf_143_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_144_clock (.I(clknet_5_24_0_clock),
    .Z(clknet_leaf_144_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_145_clock (.I(clknet_5_24_0_clock),
    .Z(clknet_leaf_145_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_146_clock (.I(clknet_5_24_0_clock),
    .Z(clknet_leaf_146_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_147_clock (.I(clknet_5_24_0_clock),
    .Z(clknet_leaf_147_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_148_clock (.I(clknet_5_24_0_clock),
    .Z(clknet_leaf_148_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_149_clock (.I(clknet_5_24_0_clock),
    .Z(clknet_leaf_149_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_150_clock (.I(clknet_5_25_0_clock),
    .Z(clknet_leaf_150_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_151_clock (.I(clknet_5_25_0_clock),
    .Z(clknet_leaf_151_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_152_clock (.I(clknet_5_25_0_clock),
    .Z(clknet_leaf_152_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_153_clock (.I(clknet_5_25_0_clock),
    .Z(clknet_leaf_153_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_154_clock (.I(clknet_5_27_0_clock),
    .Z(clknet_leaf_154_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_155_clock (.I(clknet_5_27_0_clock),
    .Z(clknet_leaf_155_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_156_clock (.I(clknet_5_26_0_clock),
    .Z(clknet_leaf_156_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_157_clock (.I(clknet_5_26_0_clock),
    .Z(clknet_leaf_157_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_158_clock (.I(clknet_5_26_0_clock),
    .Z(clknet_leaf_158_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_159_clock (.I(clknet_5_26_0_clock),
    .Z(clknet_leaf_159_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_160_clock (.I(clknet_5_26_0_clock),
    .Z(clknet_leaf_160_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_161_clock (.I(clknet_5_26_0_clock),
    .Z(clknet_leaf_161_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_162_clock (.I(clknet_5_26_0_clock),
    .Z(clknet_leaf_162_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_163_clock (.I(clknet_5_26_0_clock),
    .Z(clknet_leaf_163_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_164_clock (.I(clknet_5_26_0_clock),
    .Z(clknet_leaf_164_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_165_clock (.I(clknet_5_26_0_clock),
    .Z(clknet_leaf_165_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_166_clock (.I(clknet_5_26_0_clock),
    .Z(clknet_leaf_166_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_167_clock (.I(clknet_5_26_0_clock),
    .Z(clknet_leaf_167_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_168_clock (.I(clknet_5_27_0_clock),
    .Z(clknet_leaf_168_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_169_clock (.I(clknet_5_27_0_clock),
    .Z(clknet_leaf_169_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_170_clock (.I(clknet_5_27_0_clock),
    .Z(clknet_leaf_170_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_171_clock (.I(clknet_5_27_0_clock),
    .Z(clknet_leaf_171_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_172_clock (.I(clknet_5_27_0_clock),
    .Z(clknet_leaf_172_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_173_clock (.I(clknet_5_27_0_clock),
    .Z(clknet_leaf_173_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_174_clock (.I(clknet_5_27_0_clock),
    .Z(clknet_leaf_174_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_175_clock (.I(clknet_5_27_0_clock),
    .Z(clknet_leaf_175_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_177_clock (.I(clknet_5_27_0_clock),
    .Z(clknet_leaf_177_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_178_clock (.I(clknet_5_30_0_clock),
    .Z(clknet_leaf_178_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_179_clock (.I(clknet_5_30_0_clock),
    .Z(clknet_leaf_179_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_180_clock (.I(clknet_5_30_0_clock),
    .Z(clknet_leaf_180_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_181_clock (.I(clknet_5_30_0_clock),
    .Z(clknet_leaf_181_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_182_clock (.I(clknet_5_27_0_clock),
    .Z(clknet_leaf_182_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_183_clock (.I(clknet_5_30_0_clock),
    .Z(clknet_leaf_183_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_184_clock (.I(clknet_5_27_0_clock),
    .Z(clknet_leaf_184_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_185_clock (.I(clknet_5_30_0_clock),
    .Z(clknet_leaf_185_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_186_clock (.I(clknet_5_31_0_clock),
    .Z(clknet_leaf_186_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_187_clock (.I(clknet_5_31_0_clock),
    .Z(clknet_leaf_187_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_188_clock (.I(clknet_5_31_0_clock),
    .Z(clknet_leaf_188_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_189_clock (.I(clknet_5_31_0_clock),
    .Z(clknet_leaf_189_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_190_clock (.I(clknet_5_31_0_clock),
    .Z(clknet_leaf_190_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_191_clock (.I(clknet_5_31_0_clock),
    .Z(clknet_leaf_191_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_192_clock (.I(clknet_5_31_0_clock),
    .Z(clknet_leaf_192_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_193_clock (.I(clknet_5_31_0_clock),
    .Z(clknet_leaf_193_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_194_clock (.I(clknet_5_31_0_clock),
    .Z(clknet_leaf_194_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_195_clock (.I(clknet_5_31_0_clock),
    .Z(clknet_leaf_195_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_196_clock (.I(clknet_5_31_0_clock),
    .Z(clknet_leaf_196_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_197_clock (.I(clknet_5_30_0_clock),
    .Z(clknet_leaf_197_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_198_clock (.I(clknet_5_30_0_clock),
    .Z(clknet_leaf_198_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_199_clock (.I(clknet_5_28_0_clock),
    .Z(clknet_leaf_199_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_200_clock (.I(clknet_5_28_0_clock),
    .Z(clknet_leaf_200_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_201_clock (.I(clknet_5_28_0_clock),
    .Z(clknet_leaf_201_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_202_clock (.I(clknet_5_29_0_clock),
    .Z(clknet_leaf_202_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_203_clock (.I(clknet_5_29_0_clock),
    .Z(clknet_leaf_203_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_204_clock (.I(clknet_5_29_0_clock),
    .Z(clknet_leaf_204_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_205_clock (.I(clknet_5_29_0_clock),
    .Z(clknet_leaf_205_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_206_clock (.I(clknet_5_29_0_clock),
    .Z(clknet_leaf_206_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_207_clock (.I(clknet_5_29_0_clock),
    .Z(clknet_leaf_207_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_208_clock (.I(clknet_5_29_0_clock),
    .Z(clknet_leaf_208_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_209_clock (.I(clknet_5_29_0_clock),
    .Z(clknet_leaf_209_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_210_clock (.I(clknet_5_29_0_clock),
    .Z(clknet_leaf_210_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_211_clock (.I(clknet_5_29_0_clock),
    .Z(clknet_leaf_211_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_212_clock (.I(clknet_5_29_0_clock),
    .Z(clknet_leaf_212_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_213_clock (.I(clknet_5_29_0_clock),
    .Z(clknet_leaf_213_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_214_clock (.I(clknet_5_28_0_clock),
    .Z(clknet_leaf_214_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_215_clock (.I(clknet_5_28_0_clock),
    .Z(clknet_leaf_215_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_216_clock (.I(clknet_5_28_0_clock),
    .Z(clknet_leaf_216_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_217_clock (.I(clknet_5_28_0_clock),
    .Z(clknet_leaf_217_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_218_clock (.I(clknet_5_28_0_clock),
    .Z(clknet_leaf_218_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_219_clock (.I(clknet_5_28_0_clock),
    .Z(clknet_leaf_219_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_220_clock (.I(clknet_5_28_0_clock),
    .Z(clknet_leaf_220_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_221_clock (.I(clknet_5_28_0_clock),
    .Z(clknet_leaf_221_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_222_clock (.I(clknet_5_28_0_clock),
    .Z(clknet_leaf_222_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_223_clock (.I(clknet_5_25_0_clock),
    .Z(clknet_leaf_223_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_224_clock (.I(clknet_5_25_0_clock),
    .Z(clknet_leaf_224_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_225_clock (.I(clknet_5_25_0_clock),
    .Z(clknet_leaf_225_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_226_clock (.I(clknet_5_25_0_clock),
    .Z(clknet_leaf_226_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_227_clock (.I(clknet_5_25_0_clock),
    .Z(clknet_leaf_227_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_228_clock (.I(clknet_5_25_0_clock),
    .Z(clknet_leaf_228_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_229_clock (.I(clknet_5_25_0_clock),
    .Z(clknet_leaf_229_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_230_clock (.I(clknet_5_24_0_clock),
    .Z(clknet_leaf_230_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_231_clock (.I(clknet_5_24_0_clock),
    .Z(clknet_leaf_231_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_232_clock (.I(clknet_5_24_0_clock),
    .Z(clknet_leaf_232_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_233_clock (.I(clknet_5_18_0_clock),
    .Z(clknet_leaf_233_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_234_clock (.I(clknet_5_18_0_clock),
    .Z(clknet_leaf_234_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_235_clock (.I(clknet_5_18_0_clock),
    .Z(clknet_leaf_235_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_236_clock (.I(clknet_5_19_0_clock),
    .Z(clknet_leaf_236_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_237_clock (.I(clknet_5_19_0_clock),
    .Z(clknet_leaf_237_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_238_clock (.I(clknet_5_19_0_clock),
    .Z(clknet_leaf_238_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_239_clock (.I(clknet_5_19_0_clock),
    .Z(clknet_leaf_239_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_240_clock (.I(clknet_5_19_0_clock),
    .Z(clknet_leaf_240_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_241_clock (.I(clknet_5_19_0_clock),
    .Z(clknet_leaf_241_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_242_clock (.I(clknet_5_19_0_clock),
    .Z(clknet_leaf_242_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_243_clock (.I(clknet_5_19_0_clock),
    .Z(clknet_leaf_243_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_244_clock (.I(clknet_5_19_0_clock),
    .Z(clknet_leaf_244_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_245_clock (.I(clknet_5_22_0_clock),
    .Z(clknet_leaf_245_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_246_clock (.I(clknet_5_22_0_clock),
    .Z(clknet_leaf_246_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_248_clock (.I(clknet_5_22_0_clock),
    .Z(clknet_leaf_248_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_249_clock (.I(clknet_5_22_0_clock),
    .Z(clknet_leaf_249_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_250_clock (.I(clknet_5_22_0_clock),
    .Z(clknet_leaf_250_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_251_clock (.I(clknet_5_22_0_clock),
    .Z(clknet_leaf_251_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_252_clock (.I(clknet_5_22_0_clock),
    .Z(clknet_leaf_252_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_253_clock (.I(clknet_5_22_0_clock),
    .Z(clknet_leaf_253_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_254_clock (.I(clknet_5_23_0_clock),
    .Z(clknet_leaf_254_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_255_clock (.I(clknet_5_23_0_clock),
    .Z(clknet_leaf_255_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_256_clock (.I(clknet_5_23_0_clock),
    .Z(clknet_leaf_256_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_257_clock (.I(clknet_5_23_0_clock),
    .Z(clknet_leaf_257_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_258_clock (.I(clknet_5_23_0_clock),
    .Z(clknet_leaf_258_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_259_clock (.I(clknet_5_23_0_clock),
    .Z(clknet_leaf_259_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_260_clock (.I(clknet_5_23_0_clock),
    .Z(clknet_leaf_260_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_261_clock (.I(clknet_5_23_0_clock),
    .Z(clknet_leaf_261_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_262_clock (.I(clknet_5_23_0_clock),
    .Z(clknet_leaf_262_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_263_clock (.I(clknet_5_23_0_clock),
    .Z(clknet_leaf_263_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_264_clock (.I(clknet_5_23_0_clock),
    .Z(clknet_leaf_264_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_265_clock (.I(clknet_5_23_0_clock),
    .Z(clknet_leaf_265_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_266_clock (.I(clknet_5_23_0_clock),
    .Z(clknet_leaf_266_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_267_clock (.I(clknet_5_22_0_clock),
    .Z(clknet_leaf_267_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_268_clock (.I(clknet_5_22_0_clock),
    .Z(clknet_leaf_268_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_269_clock (.I(clknet_5_22_0_clock),
    .Z(clknet_leaf_269_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_270_clock (.I(clknet_5_20_0_clock),
    .Z(clknet_leaf_270_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_271_clock (.I(clknet_5_20_0_clock),
    .Z(clknet_leaf_271_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_272_clock (.I(clknet_5_20_0_clock),
    .Z(clknet_leaf_272_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_273_clock (.I(clknet_5_21_0_clock),
    .Z(clknet_leaf_273_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_274_clock (.I(clknet_5_21_0_clock),
    .Z(clknet_leaf_274_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_275_clock (.I(clknet_5_21_0_clock),
    .Z(clknet_leaf_275_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_276_clock (.I(clknet_5_21_0_clock),
    .Z(clknet_leaf_276_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_277_clock (.I(clknet_5_21_0_clock),
    .Z(clknet_leaf_277_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_278_clock (.I(clknet_5_21_0_clock),
    .Z(clknet_leaf_278_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_279_clock (.I(clknet_5_21_0_clock),
    .Z(clknet_leaf_279_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_280_clock (.I(clknet_5_21_0_clock),
    .Z(clknet_leaf_280_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_281_clock (.I(clknet_5_21_0_clock),
    .Z(clknet_leaf_281_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_282_clock (.I(clknet_5_21_0_clock),
    .Z(clknet_leaf_282_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_283_clock (.I(clknet_5_21_0_clock),
    .Z(clknet_leaf_283_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_284_clock (.I(clknet_5_21_0_clock),
    .Z(clknet_leaf_284_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_285_clock (.I(clknet_5_20_0_clock),
    .Z(clknet_leaf_285_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_286_clock (.I(clknet_5_20_0_clock),
    .Z(clknet_leaf_286_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_287_clock (.I(clknet_5_20_0_clock),
    .Z(clknet_leaf_287_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_288_clock (.I(clknet_5_20_0_clock),
    .Z(clknet_leaf_288_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_289_clock (.I(clknet_5_20_0_clock),
    .Z(clknet_leaf_289_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_290_clock (.I(clknet_5_20_0_clock),
    .Z(clknet_leaf_290_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_291_clock (.I(clknet_5_20_0_clock),
    .Z(clknet_leaf_291_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_292_clock (.I(clknet_5_20_0_clock),
    .Z(clknet_leaf_292_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_293_clock (.I(clknet_5_20_0_clock),
    .Z(clknet_leaf_293_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_294_clock (.I(clknet_5_20_0_clock),
    .Z(clknet_leaf_294_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_295_clock (.I(clknet_5_17_0_clock),
    .Z(clknet_leaf_295_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_296_clock (.I(clknet_5_17_0_clock),
    .Z(clknet_leaf_296_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_297_clock (.I(clknet_5_17_0_clock),
    .Z(clknet_leaf_297_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_298_clock (.I(clknet_5_17_0_clock),
    .Z(clknet_leaf_298_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_299_clock (.I(clknet_5_17_0_clock),
    .Z(clknet_leaf_299_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_300_clock (.I(clknet_5_17_0_clock),
    .Z(clknet_leaf_300_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_301_clock (.I(clknet_5_16_0_clock),
    .Z(clknet_leaf_301_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_302_clock (.I(clknet_5_16_0_clock),
    .Z(clknet_leaf_302_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_303_clock (.I(clknet_5_16_0_clock),
    .Z(clknet_leaf_303_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_304_clock (.I(clknet_5_16_0_clock),
    .Z(clknet_leaf_304_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_305_clock (.I(clknet_5_16_0_clock),
    .Z(clknet_leaf_305_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_306_clock (.I(clknet_5_16_0_clock),
    .Z(clknet_leaf_306_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_307_clock (.I(clknet_5_16_0_clock),
    .Z(clknet_leaf_307_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_309_clock (.I(clknet_5_16_0_clock),
    .Z(clknet_leaf_309_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_310_clock (.I(clknet_5_17_0_clock),
    .Z(clknet_leaf_310_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_311_clock (.I(clknet_5_17_0_clock),
    .Z(clknet_leaf_311_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_312_clock (.I(clknet_5_17_0_clock),
    .Z(clknet_leaf_312_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_313_clock (.I(clknet_5_19_0_clock),
    .Z(clknet_leaf_313_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_314_clock (.I(clknet_5_19_0_clock),
    .Z(clknet_leaf_314_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_315_clock (.I(clknet_5_18_0_clock),
    .Z(clknet_leaf_315_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_316_clock (.I(clknet_5_18_0_clock),
    .Z(clknet_leaf_316_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_317_clock (.I(clknet_5_18_0_clock),
    .Z(clknet_leaf_317_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_318_clock (.I(clknet_5_18_0_clock),
    .Z(clknet_leaf_318_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_319_clock (.I(clknet_5_18_0_clock),
    .Z(clknet_leaf_319_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_320_clock (.I(clknet_5_18_0_clock),
    .Z(clknet_leaf_320_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_321_clock (.I(clknet_5_18_0_clock),
    .Z(clknet_leaf_321_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_322_clock (.I(clknet_5_18_0_clock),
    .Z(clknet_leaf_322_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_323_clock (.I(clknet_5_18_0_clock),
    .Z(clknet_leaf_323_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_324_clock (.I(clknet_5_7_0_clock),
    .Z(clknet_leaf_324_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_325_clock (.I(clknet_5_7_0_clock),
    .Z(clknet_leaf_325_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_326_clock (.I(clknet_5_7_0_clock),
    .Z(clknet_leaf_326_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_327_clock (.I(clknet_5_7_0_clock),
    .Z(clknet_leaf_327_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_328_clock (.I(clknet_5_7_0_clock),
    .Z(clknet_leaf_328_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_329_clock (.I(clknet_5_7_0_clock),
    .Z(clknet_leaf_329_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_330_clock (.I(clknet_5_7_0_clock),
    .Z(clknet_leaf_330_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_331_clock (.I(clknet_5_7_0_clock),
    .Z(clknet_leaf_331_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_332_clock (.I(clknet_5_7_0_clock),
    .Z(clknet_leaf_332_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_333_clock (.I(clknet_5_6_0_clock),
    .Z(clknet_leaf_333_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_334_clock (.I(clknet_5_6_0_clock),
    .Z(clknet_leaf_334_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_335_clock (.I(clknet_5_5_0_clock),
    .Z(clknet_leaf_335_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_336_clock (.I(clknet_5_4_0_clock),
    .Z(clknet_leaf_336_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_337_clock (.I(clknet_5_4_0_clock),
    .Z(clknet_leaf_337_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_338_clock (.I(clknet_5_5_0_clock),
    .Z(clknet_leaf_338_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_340_clock (.I(clknet_5_5_0_clock),
    .Z(clknet_leaf_340_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_341_clock (.I(clknet_5_5_0_clock),
    .Z(clknet_leaf_341_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_342_clock (.I(clknet_5_5_0_clock),
    .Z(clknet_leaf_342_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_343_clock (.I(clknet_5_5_0_clock),
    .Z(clknet_leaf_343_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_344_clock (.I(clknet_5_5_0_clock),
    .Z(clknet_leaf_344_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_345_clock (.I(clknet_5_5_0_clock),
    .Z(clknet_leaf_345_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_346_clock (.I(clknet_5_4_0_clock),
    .Z(clknet_leaf_346_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_347_clock (.I(clknet_5_4_0_clock),
    .Z(clknet_leaf_347_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_348_clock (.I(clknet_5_4_0_clock),
    .Z(clknet_leaf_348_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_349_clock (.I(clknet_5_4_0_clock),
    .Z(clknet_leaf_349_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_350_clock (.I(clknet_5_4_0_clock),
    .Z(clknet_leaf_350_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_352_clock (.I(clknet_5_1_0_clock),
    .Z(clknet_leaf_352_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_353_clock (.I(clknet_5_1_0_clock),
    .Z(clknet_leaf_353_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_354_clock (.I(clknet_5_1_0_clock),
    .Z(clknet_leaf_354_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_355_clock (.I(clknet_5_1_0_clock),
    .Z(clknet_leaf_355_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_356_clock (.I(clknet_5_1_0_clock),
    .Z(clknet_leaf_356_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_357_clock (.I(clknet_5_1_0_clock),
    .Z(clknet_leaf_357_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_358_clock (.I(clknet_5_1_0_clock),
    .Z(clknet_leaf_358_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_359_clock (.I(clknet_5_1_0_clock),
    .Z(clknet_leaf_359_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_360_clock (.I(clknet_5_0_0_clock),
    .Z(clknet_leaf_360_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_361_clock (.I(clknet_5_0_0_clock),
    .Z(clknet_leaf_361_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_362_clock (.I(clknet_5_0_0_clock),
    .Z(clknet_leaf_362_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_363_clock (.I(clknet_5_0_0_clock),
    .Z(clknet_leaf_363_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_364_clock (.I(clknet_5_0_0_clock),
    .Z(clknet_leaf_364_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clock (.I(clock),
    .Z(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_clock (.I(clknet_0_clock),
    .Z(clknet_3_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_clock (.I(clknet_0_clock),
    .Z(clknet_3_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_clock (.I(clknet_0_clock),
    .Z(clknet_3_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_clock (.I(clknet_0_clock),
    .Z(clknet_3_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_clock (.I(clknet_0_clock),
    .Z(clknet_3_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_clock (.I(clknet_0_clock),
    .Z(clknet_3_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_clock (.I(clknet_0_clock),
    .Z(clknet_3_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_clock (.I(clknet_0_clock),
    .Z(clknet_3_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_0_0_clock (.I(clknet_3_0_0_clock),
    .Z(clknet_4_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_1_0_clock (.I(clknet_3_0_0_clock),
    .Z(clknet_4_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_2_0_clock (.I(clknet_3_1_0_clock),
    .Z(clknet_4_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_3_0_clock (.I(clknet_3_1_0_clock),
    .Z(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_4_0_clock (.I(clknet_3_2_0_clock),
    .Z(clknet_4_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_5_0_clock (.I(clknet_3_2_0_clock),
    .Z(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_6_0_clock (.I(clknet_3_3_0_clock),
    .Z(clknet_4_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_7_0_clock (.I(clknet_3_3_0_clock),
    .Z(clknet_4_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_8_0_clock (.I(clknet_3_4_0_clock),
    .Z(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_9_0_clock (.I(clknet_3_4_0_clock),
    .Z(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_10_0_clock (.I(clknet_3_5_0_clock),
    .Z(clknet_4_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_11_0_clock (.I(clknet_3_5_0_clock),
    .Z(clknet_4_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_12_0_clock (.I(clknet_3_6_0_clock),
    .Z(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_13_0_clock (.I(clknet_3_6_0_clock),
    .Z(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_14_0_clock (.I(clknet_3_7_0_clock),
    .Z(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_15_0_clock (.I(clknet_3_7_0_clock),
    .Z(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_0_0_clock (.I(clknet_4_0_0_clock),
    .Z(clknet_5_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_1_0_clock (.I(clknet_4_0_0_clock),
    .Z(clknet_5_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_2_0_clock (.I(clknet_4_1_0_clock),
    .Z(clknet_5_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_3_0_clock (.I(clknet_4_1_0_clock),
    .Z(clknet_5_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_4_0_clock (.I(clknet_4_2_0_clock),
    .Z(clknet_5_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_5_0_clock (.I(clknet_4_2_0_clock),
    .Z(clknet_5_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_6_0_clock (.I(clknet_4_3_0_clock),
    .Z(clknet_5_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_7_0_clock (.I(clknet_4_3_0_clock),
    .Z(clknet_5_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_8_0_clock (.I(clknet_4_4_0_clock),
    .Z(clknet_5_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_9_0_clock (.I(clknet_4_4_0_clock),
    .Z(clknet_5_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_10_0_clock (.I(clknet_4_5_0_clock),
    .Z(clknet_5_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_11_0_clock (.I(clknet_4_5_0_clock),
    .Z(clknet_5_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_12_0_clock (.I(clknet_4_6_0_clock),
    .Z(clknet_5_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_13_0_clock (.I(clknet_4_6_0_clock),
    .Z(clknet_5_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_14_0_clock (.I(clknet_4_7_0_clock),
    .Z(clknet_5_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_15_0_clock (.I(clknet_4_7_0_clock),
    .Z(clknet_5_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_16_0_clock (.I(clknet_4_8_0_clock),
    .Z(clknet_5_16_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_17_0_clock (.I(clknet_4_8_0_clock),
    .Z(clknet_5_17_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_18_0_clock (.I(clknet_4_9_0_clock),
    .Z(clknet_5_18_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_19_0_clock (.I(clknet_4_9_0_clock),
    .Z(clknet_5_19_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_20_0_clock (.I(clknet_4_10_0_clock),
    .Z(clknet_5_20_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_21_0_clock (.I(clknet_4_10_0_clock),
    .Z(clknet_5_21_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_22_0_clock (.I(clknet_4_11_0_clock),
    .Z(clknet_5_22_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_23_0_clock (.I(clknet_4_11_0_clock),
    .Z(clknet_5_23_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_24_0_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_5_24_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_25_0_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_5_25_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_26_0_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_5_26_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_27_0_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_5_27_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_28_0_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_5_28_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_29_0_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_5_29_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_30_0_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_5_30_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_31_0_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_5_31_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clock_a (.I(clock_a),
    .Z(clknet_0_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_clock_a (.I(clknet_0_clock_a),
    .Z(clknet_2_0__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_clock_a (.I(clknet_0_clock_a),
    .Z(clknet_2_1__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_clock_a (.I(clknet_0_clock_a),
    .Z(clknet_2_2__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_clock_a (.I(clknet_0_clock_a),
    .Z(clknet_2_3__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_4 hold1 (.I(\output_active_trans.data_sync ),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12112__D (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12118__D (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06411__S (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06002__A2 (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06001__I (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05994__S (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06011__I (.I(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__I (.I(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06009__I (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__I (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__S (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06032__S (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06007__S (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06003__A2 (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__I (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__I (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06031__B2 (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06025__A1 (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06019__B2 (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__A1 (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06029__A2 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__A2 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06017__A2 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__A2 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06033__S (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06034__A2 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06035__I (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__A1 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06038__I (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__A1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__A1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06425__A1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06219__A1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__I (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06102__A1 (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06064__A1 (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06046__A1 (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__B (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06127__A1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__A3 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06046__A2 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__A1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__A1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__A1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06046__B (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06243__I (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__B (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__I (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06409__A2 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06274__B (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__A2 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__I (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__A1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06087__A1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__I (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06050__I (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__A1 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__A1 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06105__I (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06058__A2 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__A2 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__A1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06179__A1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06057__I (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__A2 (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__I (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06071__A2 (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06181__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06096__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__I (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06153__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06138__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__I (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06064__A2 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06116__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__A2 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__B1 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06223__I (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06071__B1 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06132__A2 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06090__A1 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06076__A2 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__A2 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__C1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06225__I (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06071__C1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__A1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__A3 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__A3 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06109__I (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06074__I (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06214__A2 (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__A3 (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06144__A1 (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06076__A1 (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__A2 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A1 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06082__A1 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06179__A3 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06093__I (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06089__I (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06081__I (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__A3 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__A3 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__A3 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06082__A2 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__C1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__I (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06083__B1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__A2 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__A3 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__A2 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__A2 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06247__I (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06091__A2 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__B1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__B1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__I (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A3 (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06193__A2 (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__A2 (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06090__A2 (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__A3 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__A2 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06096__A2 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06094__A1 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__A1 (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06138__A3 (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06100__I (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06094__A2 (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__A2 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__A2 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06095__I (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__A2 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__A2 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06097__I (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__A4 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__A1 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06146__A1 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__A2 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__A2 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06103__A1 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__A2 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06125__A2 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06103__A2 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06104__I (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__A1 (.I(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A1 (.I(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__A1 (.I(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06107__A2 (.I(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06265__I (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__B1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__B1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__A2 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06193__A1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__A2 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06111__A1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06156__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A2 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06116__A2 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06111__A2 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06207__A2 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06156__A2 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__A1 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__I (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06241__A2 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__A2 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06271__I (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06241__B1 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__B1 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__A2 (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06181__A2 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06146__A2 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06123__A2 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__B1 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__B1 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__I (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__B1 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__B1 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__B1 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06130__A2 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06389__A2 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A2 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06126__I (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__A2 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06163__A2 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06144__A2 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__A2 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06389__B1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__B1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06129__I (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__A3 (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06168__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06163__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06132__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__A2 (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A2 (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06133__I (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06176__A2 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06168__A2 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__A1 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__C2 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__C2 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06136__I (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__C2 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__C2 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06139__I (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__B1 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__B1 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06224__B1 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06140__C2 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__A4 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06377__C2 (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__C2 (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__I (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06344__A2 (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__A2 (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__A2 (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__C2 (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__A2 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__A2 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__I (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06277__B1 (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__B1 (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__I (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__C1 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__C1 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06154__I (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06162__A2 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__I (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06191__A2 (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__A1 (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__A2 (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__B1 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__B1 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06160__I (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06218__A2 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06400__A2 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06365__A2 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06164__I (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06400__B1 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06365__B1 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06166__I (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06406__A2 (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__A2 (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06169__I (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06336__A2 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__A2 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06238__A2 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__A2 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__A2 (.I(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__A2 (.I(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06179__A2 (.I(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06171__I (.I(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__B2 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06214__A1 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06191__A3 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__A1 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06406__B1 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__B1 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06173__I (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06336__B1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__B1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06238__B1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__B1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__A2 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__A2 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06175__I (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__B1 (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__B1 (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06177__I (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06189__A1 (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06402__A2 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06367__A2 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06180__I (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06402__B1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06367__B1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06182__I (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__B1 (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06296__B1 (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__B1 (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__B1 (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__A2 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06369__A2 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06185__I (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__B1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06369__B1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__I (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06330__A2 (.I(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__B1 (.I(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06192__I (.I(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__A2 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__A2 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__A2 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__A2 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06330__B1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__C2 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06194__I (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__B1 (.I(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__B1 (.I(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__B1 (.I(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__B1 (.I(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__A2 (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06326__A2 (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06196__I (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__B1 (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06326__B1 (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06198__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06360__B1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06289__B1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06257__C1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06199__B1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06396__A2 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06327__A2 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__I (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06396__B1 (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06327__B1 (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__I (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__A2 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__A2 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06206__I (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__B1 (.I(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__B1 (.I(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06208__I (.I(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__B1 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06291__B1 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__A2 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__B1 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__A3 (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__A2 (.I(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__A2 (.I(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06213__I (.I(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__B1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__B1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06215__I (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06218__A3 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06219__B (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07217__A1 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06221__I (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08039__A1 (.I(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06721__A1 (.I(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06431__A1 (.I(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__A1 (.I(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__B1 (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__C1 (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__B1 (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__B1 (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06353__B1 (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__A2 (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06287__B1 (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06229__B1 (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__B1 (.I(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06237__A2 (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__A1 (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__A2 (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__A2 (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__A3 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__A3 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__A4 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06260__A3 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__A4 (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07260__A1 (.I(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__I (.I(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__A1 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06757__A1 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06437__A1 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__A1 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06275__A3 (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__A1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06279__A2 (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__A2 (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__A1 (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__A3 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__C (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__A1 (.I(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__A2 (.I(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__A4 (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__B (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07304__A1 (.I(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__I (.I(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__A1 (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__A1 (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__A1 (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__A1 (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A2 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06338__A1 (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06322__A2 (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06324__A4 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06338__A3 (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06330__C (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06337__A2 (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__A2 (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06338__A4 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__B (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07391__A1 (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__I (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__A1 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__A1 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__A1 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06374__A1 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06345__A2 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06373__A1 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06350__A2 (.I(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06373__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__C (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06373__A3 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__C (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06372__A1 (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06372__A2 (.I(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06373__A4 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06374__B (.I(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07454__A1 (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__I (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__A1 (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06858__A1 (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06449__A1 (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06409__A1 (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__A2 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06408__A1 (.I(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__A2 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06408__A2 (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06394__A2 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__C (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06408__A3 (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__A1 (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06408__A4 (.I(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06409__B (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06497__C (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__I (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__A1 (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__A1 (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__I (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__A2 (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06473__I (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__I (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06419__I (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06413__I (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__I (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__I (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__C (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__I (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__A2 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06437__A2 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06431__A2 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06425__A2 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06497__A2 (.I(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06491__A2 (.I(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06487__A2 (.I(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__A2 (.I(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__I (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__I (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__I (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__I (.I(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__I (.I(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__I (.I(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__I (.I(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06498__A2 (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__A2 (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__A2 (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__A2 (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06496__A2 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__I (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06446__I (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__I (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06482__A2 (.I(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06467__A2 (.I(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__B1 (.I(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__B1 (.I(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06463__A2 (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06445__A2 (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__A2 (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06433__A2 (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06490__A2 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__A2 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__B1 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06436__B1 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__C (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__C (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__C (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06436__C (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06437__B2 (.I(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__B2 (.I(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06460__A2 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__A2 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06449__A2 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__A2 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__A2 (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__A2 (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06455__A2 (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__A2 (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__B1 (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__B1 (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__B1 (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__B1 (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06449__B2 (.I(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__A1 (.I(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A1 (.I(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__A1 (.I(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__B1 (.I(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__B1 (.I(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__B1 (.I(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__B1 (.I(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06455__B1 (.I(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A1 (.I(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A1 (.I(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06460__A1 (.I(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06460__B1 (.I(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__A1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__A1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06465__A1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__A2 (.I(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__A2 (.I(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__A2 (.I(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06465__A2 (.I(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08071__A1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07691__A1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__A1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__A2 (.I(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__A2 (.I(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__A2 (.I(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__A2 (.I(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__A1 (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__A1 (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__A1 (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06487__C (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__C (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__C (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__C (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08077__A1 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07778__A1 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__A1 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__A1 (.I(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__A1 (.I(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__A1 (.I(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06498__B1 (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__A2 (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__A2 (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__A2 (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__B2 (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A1 (.I(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07908__A1 (.I(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__A1 (.I(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__A1 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__A1 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__A1 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__A1 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__A1 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06498__B2 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11912__A1 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06496__A1 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06648__A1 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06616__A1 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06603__A1 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06508__B (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__B (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06698__B (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__I (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__A2 (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__B (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06721__A2 (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__I (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06672__A2 (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__A2 (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__A1 (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__I (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A2 (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06631__A1 (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06557__A2 (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__A1 (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__A2 (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06629__A2 (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06616__A2 (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__A2 (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__A1 (.I(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06572__I (.I(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__I (.I(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__I (.I(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__A1 (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06613__A1 (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__A1 (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__A1 (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__A2 (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__A2 (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__A2 (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06779__B1 (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__B1 (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__I (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06606__A2 (.I(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__A1 (.I(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06553__A1 (.I(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06534__A1 (.I(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A2 (.I(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__A2 (.I(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06534__A2 (.I(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__B1 (.I(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__C1 (.I(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__I (.I(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__A1 (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__I (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__I (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__I (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__A1 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06601__A1 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__A1 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__A1 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A2 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06540__I (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06615__A1 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__A2 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__A2 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__A2 (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06780__A2 (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06545__I (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__A2 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06728__A2 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__A2 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__A2 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__A1 (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__A1 (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06565__A1 (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__A1 (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__A2 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06601__A2 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__A2 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__B1 (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__B1 (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__I (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__A2 (.I(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06561__A2 (.I(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__A1 (.I(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06552__A2 (.I(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06624__A2 (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__A2 (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06553__A2 (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__C2 (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__C2 (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06554__I (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06564__A2 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__A2 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06565__A2 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06557__A1 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06833__A2 (.I(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06779__A2 (.I(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__I (.I(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06651__A2 (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A1 (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06596__A1 (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06560__I (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A2 (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06708__I (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__B1 (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__A1 (.I(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__A2 (.I(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06648__A2 (.I(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__A2 (.I(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__A1 (.I(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__A1 (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06615__A2 (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__A2 (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__A2 (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__A2 (.I(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__A1 (.I(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06574__A2 (.I(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06589__A2 (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__A2 (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__A2 (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__I (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__B1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__B1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06583__I (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__A2 (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__A2 (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__A2 (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__A2 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__A2 (.I(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__A2 (.I(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06591__I (.I(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__A2 (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__A2 (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__A2 (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__B1 (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__B1 (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__I (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06613__A2 (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06606__A1 (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06603__A2 (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06596__A2 (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06777__A2 (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__C2 (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06597__I (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__A2 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__A2 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__I (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__B1 (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__B1 (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__I (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__B1 (.I(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__C2 (.I(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__I (.I(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06841__C2 (.I(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06739__B1 (.I(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__C2 (.I(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__C2 (.I(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__A2 (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06777__B1 (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06607__I (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__C1 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06739__A2 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06705__C1 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06610__A2 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__C2 (.I(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06774__A2 (.I(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06609__I (.I(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__A2 (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__A2 (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__I (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__B1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__B1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06614__I (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06835__A2 (.I(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__I (.I(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__A2 (.I(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__A2 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06701__I (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__A2 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__A1 (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A2 (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06620__A2 (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__B1 (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06693__I (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__B1 (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__A1 (.I(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__A1 (.I(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__A1 (.I(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06624__A1 (.I(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__C (.I(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__A4 (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__A3 (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__A2 (.I(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__C2 (.I(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06630__I (.I(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__B1 (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__B1 (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__I (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__A2 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__A2 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__I (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__B1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06787__B1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__I (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06672__A1 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__A2 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06641__A2 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__I (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__A2 (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__A2 (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06743__I (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__C1 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__B1 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__A2 (.I(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__A2 (.I(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06644__I (.I(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__B1 (.I(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__B1 (.I(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06646__I (.I(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__A2 (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06714__I (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__A2 (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__B1 (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__I (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__B1 (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06846__A2 (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06712__I (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__A2 (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06846__B1 (.I(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06716__I (.I(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__B1 (.I(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06677__A3 (.I(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__A2 (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__A2 (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06657__I (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__A2 (.I(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__A2 (.I(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__A2 (.I(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__A2 (.I(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__B1 (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__B1 (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06659__I (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__B1 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__B1 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__B1 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__B1 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06851__A2 (.I(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__A2 (.I(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__I (.I(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06851__B1 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__B1 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__I (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06852__A2 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__A2 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06666__I (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06852__B1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__B1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06668__I (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06675__A2 (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06853__A2 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__A2 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06671__I (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__A2 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06787__A2 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06686__A2 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__A2 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06853__B1 (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__B1 (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06673__I (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__A4 (.I(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__B (.I(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__A2 (.I(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06721__B1 (.I(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06695__A1 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__C2 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__A2 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__A2 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__C2 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06695__A4 (.I(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__A1 (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__A1 (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__A2 (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__A3 (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__A3 (.I(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06719__A3 (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06719__A4 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__A4 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06721__B2 (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__A2 (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__A1 (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__A2 (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__A2 (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__A1 (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__A1 (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__A3 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__A1 (.I(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__C (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__A2 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__A3 (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__A4 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06757__B (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06761__A2 (.I(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__B1 (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__A1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__A2 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__A3 (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06773__A2 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06789__A1 (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06778__A2 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06789__A2 (.I(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__A2 (.I(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06789__A4 (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__B2 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06804__A1 (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06800__A1 (.I(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06804__A2 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06804__A3 (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06804__A4 (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__A1 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06809__A3 (.I(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__A2 (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__C (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__A3 (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__A3 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__B (.I(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06829__A3 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06834__A2 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__A2 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__C (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__A3 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__A2 (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__A4 (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06858__B (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__A2 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__A2 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__A1 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__A1 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__A1 (.I(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__A1 (.I(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__A1 (.I(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06866__A1 (.I(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__A3 (.I(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__A3 (.I(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06866__A2 (.I(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__I (.I(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06933__I (.I(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__I (.I(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07072__I (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07068__I (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__I (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__A1 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06961__A1 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__A1 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__I (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06944__A2 (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__A2 (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__A2 (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__I (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__A2 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06930__A1 (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__A1 (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__A1 (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__A1 (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06908__A3 (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__B (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__I (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__A2 (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__A2 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__A3 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__I (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06879__I (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__B (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07506__I (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07269__I (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__I (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__B (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__B (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__B (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__I (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__I (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__I (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07305__I (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__I (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07304__A2 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07260__A2 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07217__A2 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__A2 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06990__I (.I(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__I (.I(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__I (.I(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__I (.I(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07089__I (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06919__I (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06915__I (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06885__I (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07147__C (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07142__C (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06981__C (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__A1 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06908__A1 (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__A1 (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__I (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07058__I (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06959__I (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06920__I (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__I (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07137__A2 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__A2 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07069__A2 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__A2 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06953__I (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__I (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06930__A2 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__A2 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06922__I (.I(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06899__I (.I(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__A2 (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__A2 (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07028__A2 (.I(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07005__A3 (.I(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06984__A3 (.I(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__A2 (.I(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__A3 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__A3 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__A3 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__A3 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07139__A4 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06995__B (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__A4 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07781__I (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07544__I (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__I (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__I (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06987__I (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__I (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06928__I (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__I (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06988__I (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06940__I (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__I (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__I (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__A2 (.I(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A2 (.I(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06955__A2 (.I(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06914__A2 (.I(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07028__A3 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__A3 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06932__A3 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06914__A3 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__B (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07023__A4 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A4 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06916__B (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__C (.I(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__C (.I(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07041__A1 (.I(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06916__C (.I(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__I (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__I (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07308__I (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06917__I (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__A1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06985__C (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__A1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06926__A1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__A1 (.I(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06984__A2 (.I(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06955__A1 (.I(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__A1 (.I(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06942__I (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06924__I (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__A2 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__A2 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06932__A2 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__A2 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07132__B (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__B (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A4 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06926__A4 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__I (.I(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07547__I (.I(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07310__I (.I(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__I (.I(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__A1 (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__A1 (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06972__I (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__A1 (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__A2 (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__A2 (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06973__I (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__A2 (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06932__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07069__A4 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__A4 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__B (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__B (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__I (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__I (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__I (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__I (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07051__A1 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A1 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A1 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__C (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07785__I (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__I (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__I (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06936__I (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07098__I (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__I (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06979__I (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06939__I (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07099__I (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07088__I (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__I (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__I (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06944__A1 (.I(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06961__A2 (.I(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06945__A2 (.I(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A3 (.I(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06974__A3 (.I(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06955__A3 (.I(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06946__A3 (.I(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07090__B (.I(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07062__A4 (.I(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A4 (.I(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06948__B (.I(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__C (.I(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07102__C (.I(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07062__A1 (.I(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06948__C (.I(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07787__I (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__I (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__I (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__I (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__A2 (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__A2 (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07160__A2 (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__A2 (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07043__A1 (.I(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__A1 (.I(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A1 (.I(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06956__A1 (.I(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__I (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__I (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__I (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__I (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__I (.I(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07013__I (.I(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__I (.I(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06954__I (.I(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07149__A3 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07051__A3 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A3 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06956__A3 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__B (.I(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__A4 (.I(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07000__B (.I(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06956__A4 (.I(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__I (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__I (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__I (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06957__I (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__B1 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__B1 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07160__B1 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__B1 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07073__A1 (.I(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07005__A1 (.I(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06984__A1 (.I(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06963__A1 (.I(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07028__A1 (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07005__A2 (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06974__A1 (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06963__A2 (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__B (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07079__A4 (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06981__B (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__A4 (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07629__I (.I(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07392__I (.I(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07155__I (.I(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06965__I (.I(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__A2 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__A2 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__A2 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06970__A2 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07043__A2 (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A2 (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__A2 (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A2 (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07043__A3 (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A3 (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__A3 (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A3 (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07630__I (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07393__I (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07156__I (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06969__I (.I(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__B1 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__B1 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__B1 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06970__B1 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__A4 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07057__A1 (.I(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A1 (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__A1 (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07000__A1 (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A1 (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A2 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__A2 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07000__A2 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A2 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07144__A4 (.I(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07107__B (.I(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07081__A4 (.I(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__B (.I(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__A1 (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__C (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__A1 (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06976__I (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__C (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07060__A1 (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07000__C (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__C (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__I (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07554__I (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07317__I (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06978__I (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__A2 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__A2 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07162__A2 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A2 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__I (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07555__I (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07318__I (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__I (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__B1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__B1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07162__B1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__B1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07111__B (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07051__A4 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__A4 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06985__B (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__I (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07557__I (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07320__I (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__I (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__A1 (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__A1 (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__A1 (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__A1 (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__A2 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__A2 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__A2 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__A2 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07137__A4 (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__B (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07031__A4 (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__B (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__I (.I(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__I (.I(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__I (.I(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06992__I (.I(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07267__B1 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07224__B1 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07163__B1 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__B1 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07003__A2 (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07139__A1 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07107__C (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07081__A1 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06995__C (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07797__I (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__I (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__I (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06996__I (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07225__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__I (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07561__I (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07324__I (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__I (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__B1 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07225__B1 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__B1 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__B1 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__I (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__I (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07326__I (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__I (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__A2 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__A2 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__A2 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__A2 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07057__A2 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__C (.I(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07123__C (.I(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07023__A1 (.I(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07006__A1 (.I(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07147__B (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07123__B (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07060__A4 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07006__A4 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07805__I (.I(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07568__I (.I(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__I (.I(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__I (.I(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__A2 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__A2 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__A2 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__A2 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__C (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07031__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__I (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07569__I (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07332__I (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07010__I (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__B1 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__B1 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__B1 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__B1 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07095__B (.I(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__B (.I(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07043__A4 (.I(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A4 (.I(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__I (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07571__I (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07334__I (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__I (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A2 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__A2 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07174__A2 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07022__A2 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__B (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__A4 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__B (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__A4 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07809__I (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__I (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__I (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07021__I (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07034__A2 (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07641__I (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07404__I (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__I (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07024__I (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07962__A2 (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__A2 (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__A2 (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07027__A2 (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07642__I (.I(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__I (.I(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__I (.I(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__I (.I(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07962__B1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__B1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__B1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07027__B1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07149__A4 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07142__B (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__B (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A4 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07644__I (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07407__I (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07170__I (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__I (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__A2 (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A2 (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__A2 (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__A2 (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__I (.I(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__I (.I(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07171__I (.I(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07032__I (.I(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__B1 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__B1 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__B1 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__B1 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07057__A3 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07815__I (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07578__I (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07341__I (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07036__I (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__A2 (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__A2 (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__A2 (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__A2 (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__I (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__I (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07342__I (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__I (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__B1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__B1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__B1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__B1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__B (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07066__A4 (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__B (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07041__A4 (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__I (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07413__I (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__I (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07042__I (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__A2 (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__A2 (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07881__A2 (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__A2 (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__B1 (.I(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__B1 (.I(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07881__B1 (.I(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__B1 (.I(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07653__I (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__I (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07179__I (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07047__I (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__A2 (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__A2 (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__A2 (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07050__A2 (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07654__I (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__I (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__I (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07049__I (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__B1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__B1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__B1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07050__B1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07656__I (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__I (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07182__I (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07052__I (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A2 (.I(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A2 (.I(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07883__A2 (.I(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07055__A2 (.I(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__I (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07420__I (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07183__I (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07054__I (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__B1 (.I(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__B1 (.I(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07883__B1 (.I(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07055__B1 (.I(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07057__A4 (.I(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07824__I (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__I (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07350__I (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__I (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__A2 (.I(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__A2 (.I(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__A2 (.I(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07064__A2 (.I(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__I (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__I (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07351__I (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__I (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__B1 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__B1 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__B1 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07064__B1 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07111__C (.I(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__C (.I(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__C (.I(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07066__A1 (.I(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07821__I (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__I (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__I (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07067__I (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07284__A2 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__A2 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__A2 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07071__A2 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__C (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__A1 (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__C (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07069__A1 (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__I (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07585__I (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07348__I (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07070__I (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07284__B1 (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__B1 (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__B1 (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07071__B1 (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__C (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__C (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07079__A1 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__A1 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07102__B (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__B (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__A4 (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__A4 (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07827__I (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__I (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07353__I (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07075__I (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__A2 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07242__A2 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07193__A2 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07078__A2 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__I (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__I (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__I (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07077__I (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__B1 (.I(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07242__B1 (.I(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07193__B1 (.I(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07078__B1 (.I(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__I (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__I (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07188__I (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07080__I (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__A2 (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__A2 (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07887__A2 (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07083__A2 (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__I (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__I (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07189__I (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07082__I (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__B1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__B1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07887__B1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07083__B1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07153__A1 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__I (.I(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07595__I (.I(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07358__I (.I(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07086__I (.I(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07289__A2 (.I(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__A2 (.I(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__A2 (.I(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07092__A2 (.I(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07137__A1 (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07132__C (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07095__C (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07090__C (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__I (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__I (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07359__I (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07091__I (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07289__B1 (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__B1 (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__B1 (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07092__B1 (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07669__I (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07432__I (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__I (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07094__I (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__A2 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__A2 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A2 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__A2 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07670__I (.I(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07433__I (.I(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__I (.I(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__I (.I(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__B1 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__B1 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__B1 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__B1 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__I (.I(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07598__I (.I(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07361__I (.I(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07101__I (.I(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A2 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__A2 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__A2 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07104__A2 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__I (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07599__I (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07362__I (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__I (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__B1 (.I(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__B1 (.I(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__B1 (.I(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07104__B1 (.I(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__I (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__I (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07364__I (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07106__I (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__A2 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__A2 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__A2 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__A2 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__I (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__I (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07365__I (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07108__I (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__B1 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__B1 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__B1 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__B1 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07153__A2 (.I(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__I (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__I (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__I (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07112__I (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__A2 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__A2 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A2 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07115__A2 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__I (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__I (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07370__I (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07114__I (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__B1 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__B1 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__B1 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07115__B1 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__I (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07439__I (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__I (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07117__I (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__A2 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__A2 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__A2 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07120__A2 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__I (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07440__I (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07203__I (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07119__I (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__B1 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__B1 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__B1 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07120__B1 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__I (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__I (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07372__I (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07122__I (.I(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07295__A2 (.I(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07251__A2 (.I(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__A2 (.I(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07125__A2 (.I(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07847__I (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07610__I (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07373__I (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__I (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07295__B1 (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07251__B1 (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__B1 (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07125__B1 (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07849__I (.I(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__I (.I(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07375__I (.I(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07127__I (.I(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__A2 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__A2 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__A2 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07130__A2 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__I (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07613__I (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__I (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__I (.I(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__B1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__B1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__B1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07130__B1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07153__A3 (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__I (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__I (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__I (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__I (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__A2 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__A2 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__A2 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07136__A2 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__I (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__I (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07384__I (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07135__I (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__B1 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__B1 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__B1 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07136__B1 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__I (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__I (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07380__I (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07138__I (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07299__A2 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__A2 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07212__A2 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07141__A2 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__I (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07618__I (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__I (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07140__I (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07299__B1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__B1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07212__B1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07141__B1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07860__I (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__I (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07386__I (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07143__I (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07301__A2 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07257__A2 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07214__A2 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07146__A2 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07861__I (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__I (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07387__I (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07145__I (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07301__B1 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07257__B1 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07214__B1 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07146__B1 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__I (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__I (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07209__I (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07148__I (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__A2 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A2 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__A2 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07151__A2 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__B1 (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__B1 (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__B1 (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07151__B1 (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07153__A4 (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07306__A2 (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07261__A2 (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__A2 (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__A2 (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07306__B1 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07261__B1 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__B1 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__B1 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__A1 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07166__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07329__A2 (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07272__A2 (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__A2 (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__A2 (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07329__B1 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07272__B1 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__B1 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__B1 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07330__A2 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07273__A2 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__A2 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07172__A2 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07330__B1 (.I(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07273__B1 (.I(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__B1 (.I(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07172__B1 (.I(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__A3 (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07338__A2 (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__A2 (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__A2 (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__A2 (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07338__B1 (.I(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__B1 (.I(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__B1 (.I(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__B1 (.I(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07339__A2 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__A2 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__A2 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__A2 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07339__B1 (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__B1 (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__B1 (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__B1 (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07340__A2 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__A2 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__A2 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07184__A2 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07340__B1 (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__B1 (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__B1 (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07184__B1 (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__A4 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07217__B1 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07346__A2 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07283__A2 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__A2 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07190__A2 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07346__B1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07283__B1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__B1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07190__B1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__A1 (.I(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07216__A1 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07357__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07244__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07197__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07357__B1 (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__B1 (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07244__B1 (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07197__B1 (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07216__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07368__A2 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07293__A2 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__A2 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07204__A2 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07368__B1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07293__B1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__B1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07204__B1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07216__A3 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__A2 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07298__A2 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__A2 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__A2 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__B1 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07298__B1 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__B1 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__B1 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07216__A4 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A1 (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A2 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A3 (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A4 (.I(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07260__B1 (.I(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__A1 (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__A2 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__A1 (.I(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__A2 (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__A3 (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__A4 (.I(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07282__A1 (.I(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07271__A2 (.I(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__B (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07402__B (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__B (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__B (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07282__A3 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07282__A4 (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07304__B1 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A1 (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07297__A3 (.I(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A3 (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07302__A1 (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07302__A2 (.I(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07316__A3 (.I(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07345__A1 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07328__A2 (.I(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07337__A1 (.I(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07345__A3 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07344__A4 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07345__A4 (.I(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07391__B1 (.I(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__A1 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__A2 (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__A1 (.I(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07367__A4 (.I(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__A2 (.I(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__A1 (.I(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__A4 (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__A3 (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__A4 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__A2 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__A2 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__A2 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__A2 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__B1 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__B1 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__B1 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__B1 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07424__A1 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07424__A2 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__A1 (.I(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__A2 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07510__A2 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__A2 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__A2 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__B1 (.I(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07510__B1 (.I(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__B1 (.I(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__B1 (.I(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__A3 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07424__A3 (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__A2 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__A2 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07470__A2 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__A2 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__B1 (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__B1 (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07470__B1 (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__B1 (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__A2 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__A2 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__A2 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07418__A2 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__B1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__B1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__B1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07418__B1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__B1 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__B1 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__B1 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__B1 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07424__A4 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07454__B1 (.I(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07583__A2 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A2 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__A2 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__A2 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07583__B1 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__B1 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__B1 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__B1 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07431__A2 (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__A1 (.I(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07594__A2 (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__A2 (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__A2 (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__A2 (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07594__B1 (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__B1 (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__B1 (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__B1 (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07438__A4 (.I(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__A2 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07605__A2 (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__A2 (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__A2 (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A2 (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07605__B1 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__B1 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__B1 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__B1 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07445__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__A3 (.I(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__A2 (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__A2 (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__A2 (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__A2 (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__B1 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__B1 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__B1 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__B1 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07452__A3 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__A4 (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__A1 (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A1 (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__A2 (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__A1 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__A3 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__A3 (.I(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__A4 (.I(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__B1 (.I(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07480__A2 (.I(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__A4 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A2 (.I(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A3 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07495__A3 (.I(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A4 (.I(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07502__A4 (.I(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07519__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A1 (.I(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07700__B (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07639__B (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07564__B (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__B (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07513__A1 (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07513__A3 (.I(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07519__A3 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07519__A4 (.I(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__B1 (.I(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__A2 (.I(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__A1 (.I(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__A4 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__A2 (.I(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A1 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A4 (.I(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__A3 (.I(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__A3 (.I(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__A4 (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07778__A2 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__A2 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07691__A2 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__A2 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__A2 (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A2 (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A2 (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07552__A2 (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__B1 (.I(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__B1 (.I(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__B1 (.I(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07552__B1 (.I(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A1 (.I(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07741__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07559__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07741__B1 (.I(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__B1 (.I(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__B1 (.I(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07559__B1 (.I(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07742__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07562__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07742__B1 (.I(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__B1 (.I(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__B1 (.I(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07562__B1 (.I(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__A2 (.I(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07700__A2 (.I(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07639__A2 (.I(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07564__A2 (.I(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A2 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07574__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07574__A2 (.I(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07748__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07704__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07748__B1 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07704__B1 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__B1 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__B1 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07574__A4 (.I(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A3 (.I(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__B1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__B1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__B1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__B1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__A4 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A4 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A1 (.I(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__A2 (.I(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07714__A2 (.I(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07665__A2 (.I(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__A2 (.I(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__B1 (.I(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07714__B1 (.I(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07665__B1 (.I(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__B1 (.I(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__A1 (.I(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__A2 (.I(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__A2 (.I(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__A2 (.I(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__A2 (.I(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__B1 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__B1 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__B1 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__B1 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07720__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07673__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07600__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__B1 (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07720__B1 (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07673__B1 (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07600__B1 (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__A2 (.I(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__A2 (.I(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07674__A2 (.I(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__A2 (.I(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__B1 (.I(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__B1 (.I(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07674__B1 (.I(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__B1 (.I(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__A2 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07615__A1 (.I(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__A2 (.I(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07724__A2 (.I(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__A2 (.I(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07608__A2 (.I(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__B1 (.I(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07724__B1 (.I(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__B1 (.I(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07608__B1 (.I(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__A2 (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__A2 (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07680__A2 (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__A2 (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__B1 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__B1 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07680__B1 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__B1 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__A2 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07726__A2 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__A2 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07614__A2 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__B1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07726__B1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__B1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07614__B1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__A3 (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__A2 (.I(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07729__A2 (.I(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__A2 (.I(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__A2 (.I(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__B1 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07729__B1 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__B1 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__B1 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07622__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__B1 (.I(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__B1 (.I(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__B1 (.I(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07622__B1 (.I(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__A3 (.I(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A2 (.I(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07731__A2 (.I(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07688__A2 (.I(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__A2 (.I(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__B1 (.I(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07731__B1 (.I(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07688__B1 (.I(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__B1 (.I(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__A2 (.I(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07735__A2 (.I(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__A2 (.I(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__A2 (.I(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__B1 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07735__B1 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__B1 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__B1 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07635__A2 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__A1 (.I(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__A2 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__A2 (.I(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07746__A2 (.I(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07702__A2 (.I(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__A2 (.I(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__B1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07746__B1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07702__B1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__B1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__A2 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__A2 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__A2 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__A2 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__B1 (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__B1 (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__B1 (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__B1 (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07649__A3 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__A3 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07812__A2 (.I(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__A2 (.I(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A2 (.I(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__A2 (.I(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07812__B1 (.I(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__B1 (.I(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__B1 (.I(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__B1 (.I(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__A2 (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__A2 (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07708__A2 (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07655__A2 (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__B1 (.I(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__B1 (.I(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07708__B1 (.I(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07655__B1 (.I(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07814__A2 (.I(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__A2 (.I(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__A2 (.I(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07658__A2 (.I(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07814__B1 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__B1 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__B1 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07658__B1 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__A2 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A2 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__A2 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07664__A2 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__B1 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__B1 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__B1 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07664__B1 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07668__A1 (.I(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__A1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07831__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07718__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07831__B1 (.I(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__B1 (.I(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07718__B1 (.I(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__B1 (.I(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__A2 (.I(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__A2 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07767__A2 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07723__A2 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__A2 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__B1 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07767__B1 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07723__B1 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__B1 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07682__A1 (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__A3 (.I(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07853__A2 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__A2 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__A2 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__A2 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07853__B1 (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__B1 (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__B1 (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__B1 (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__A2 (.I(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__A4 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__A2 (.I(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__A3 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__A3 (.I(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__A1 (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__A1 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__A2 (.I(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__A3 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__A4 (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__A1 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__B (.I(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__B (.I(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07801__B (.I(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__B (.I(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__A2 (.I(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__A3 (.I(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__A3 (.I(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__A1 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07777__A1 (.I(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07777__A2 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07777__A3 (.I(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__A2 (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07777__A4 (.I(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__A2 (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__A2 (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07908__A2 (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__A2 (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07790__A2 (.I(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A1 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A2 (.I(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__A2 (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A3 (.I(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A4 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__A1 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__A2 (.I(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__A3 (.I(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07864__A1 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__A4 (.I(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07864__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A1 (.I(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A3 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07864__A3 (.I(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__A2 (.I(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__A3 (.I(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07864__A4 (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__A2 (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A1 (.I(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__A2 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A2 (.I(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__A2 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A3 (.I(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A4 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__A3 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__A4 (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07901__A1 (.I(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A3 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__A2 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__A3 (.I(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A4 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__A1 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__A1 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__A2 (.I(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__A1 (.I(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__A3 (.I(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__A4 (.I(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__A1 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__A3 (.I(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__A1 (.I(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__A4 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__A2 (.I(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07944__A1 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__A3 (.I(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A2 (.I(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A3 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__A4 (.I(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__A1 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A1 (.I(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07966__A2 (.I(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A3 (.I(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A4 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07977__A1 (.I(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07977__A3 (.I(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A1 (.I(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__A4 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A2 (.I(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__A1 (.I(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__A3 (.I(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A3 (.I(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A2 (.I(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A3 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A4 (.I(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A2 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__A2 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A2 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__A2 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__B1 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__B1 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__B1 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__B1 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__A2 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__A2 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A2 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__A2 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__B1 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__B1 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__B1 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__B1 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A2 (.I(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A1 (.I(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A2 (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__B (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__A1 (.I(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__I (.I(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A1 (.I(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__A1 (.I(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__A1 (.I(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A1 (.I(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__A1 (.I(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A3 (.I(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08101__A1 (.I(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__A1 (.I(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__I (.I(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__I (.I(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__A2 (.I(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11622__A1 (.I(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11363__A1 (.I(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11104__A1 (.I(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A2 (.I(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08032__I (.I(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__I (.I(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__I (.I(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__I (.I(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__I (.I(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__I (.I(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11454__I (.I(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11195__I (.I(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__I (.I(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08031__I (.I(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11878__I1 (.I(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__I1 (.I(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__I (.I(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__A1 (.I(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__I (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__I (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__I (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__I (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11460__I (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11201__I (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__I (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08037__I (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11880__I1 (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__I1 (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__I (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__A1 (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11464__I (.I(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__I (.I(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__I (.I(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__I (.I(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11883__I1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__I1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__I (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08042__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11468__I (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__I (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__I (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__I (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11885__I1 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__I1 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__I (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08046__A1 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11472__I (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11213__I (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__I (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__I (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11887__I1 (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10811__I1 (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__I (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A1 (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11476__I (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11217__I (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08304__I (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__I (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11889__I1 (.I(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__I1 (.I(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08118__I (.I(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A1 (.I(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11892__I1 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__I1 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__I (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08059__A1 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11894__I1 (.I(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__I1 (.I(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__I (.I(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08062__A1 (.I(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08077__A2 (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__A2 (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08071__A2 (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__A2 (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11896__I1 (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10820__I1 (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__I (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__A1 (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A2 (.I(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A2 (.I(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A2 (.I(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__A2 (.I(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11898__I1 (.I(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__I1 (.I(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__I (.I(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A1 (.I(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11901__I1 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10824__I1 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08134__I (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A1 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11903__I1 (.I(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__I1 (.I(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__I (.I(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A1 (.I(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11905__I1 (.I(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__I1 (.I(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08140__I (.I(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__A1 (.I(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11907__I1 (.I(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10831__I1 (.I(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__I (.I(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__A1 (.I(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11909__I1 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10833__I1 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08147__I (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__A1 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11986__A1 (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11911__A1 (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08150__I (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08090__A1 (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__I0 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__I0 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__I0 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__I0 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08278__I (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__I (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__I (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__A3 (.I(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__A2 (.I(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__A2 (.I(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08101__A3 (.I(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__I (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__I (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__I (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__I (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__S (.I(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__S (.I(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__S (.I(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__S (.I(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__I0 (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__I0 (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__I0 (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__I0 (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__I0 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__I0 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__I0 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__I0 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__I0 (.I(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__I0 (.I(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__I0 (.I(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__I0 (.I(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08249__I0 (.I(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__I0 (.I(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__I0 (.I(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__I0 (.I(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__S (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__S (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__S (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__S (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__I0 (.I(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08209__I0 (.I(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__I0 (.I(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__I0 (.I(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__I0 (.I(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__I0 (.I(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__I0 (.I(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__I0 (.I(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__I0 (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__I0 (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__I0 (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__I0 (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__I0 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__I0 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__I0 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__I0 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__S (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__S (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__S (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__S (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__I0 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08218__I0 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__I0 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__I0 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__I0 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__I0 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08180__I0 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__I0 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__I0 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__I0 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08182__I0 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__I0 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__I0 (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__I0 (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__I0 (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__I0 (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__I0 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08227__I0 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__I0 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__I0 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__I0 (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__I0 (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__I0 (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__I0 (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08273__I0 (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__I0 (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__I0 (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__I0 (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11950__A1 (.I(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__I (.I(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08155__I (.I(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__A1 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A1 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__A1 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__I (.I(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__I (.I(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08166__I (.I(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__I (.I(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__S (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__S (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__S (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__S (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08182__S (.I(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08180__S (.I(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__S (.I(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__S (.I(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__S (.I(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__S (.I(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__S (.I(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__S (.I(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__A1 (.I(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08572__A1 (.I(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A1 (.I(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A1 (.I(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08572__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08224__I (.I(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08215__I (.I(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__I (.I(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08197__I (.I(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__S (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__S (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__S (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__S (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__S (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__S (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08209__S (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__S (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__S (.I(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__S (.I(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08218__S (.I(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__S (.I(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09321__A1 (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__A1 (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__A1 (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__A1 (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__A3 (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A3 (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__A3 (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__A3 (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__I (.I(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__I (.I(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__I (.I(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08239__I (.I(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__S (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__S (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__S (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__S (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__S (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__S (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__S (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__S (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11839__I (.I(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11776__I (.I(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11713__I (.I(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__I (.I(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__I (.I(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__I (.I(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__I (.I(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__I (.I(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08447__I0 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__I0 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__I0 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__I0 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__I (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08322__I (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08301__I (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__I (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__S (.I(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__S (.I(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__S (.I(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__S (.I(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11844__I (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11781__I (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11718__I (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08284__I (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08830__I (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__I (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08487__I (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__I (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__I0 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__I0 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__I0 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__I0 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11847__I (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11784__I (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11721__I (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__I (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08833__I (.I(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__I (.I(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__I (.I(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08290__I (.I(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08451__I0 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__I0 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__I0 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__I0 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11850__I (.I(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11787__I (.I(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11724__I (.I(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__I (.I(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__I (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__I (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__I (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08295__I (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08453__I0 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__I0 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__I0 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__I0 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11853__I (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11790__I (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11727__I (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08299__I (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__I (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__I (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__I (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__I (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__I0 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__I0 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__I0 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__I0 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__S (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__S (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__S (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__S (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11856__I (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11793__I (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11730__I (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08305__I (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__I (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__I (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__I (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__I (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__I0 (.I(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__I0 (.I(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__I0 (.I(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__I0 (.I(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10731__I (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10566__I (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__I (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08310__I (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__I (.I(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__I (.I(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__I (.I(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__I (.I(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__I0 (.I(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__I0 (.I(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__I0 (.I(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__I0 (.I(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10734__I (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10569__I (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__I (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__I (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__I (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__I (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__I (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__I (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__I0 (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08422__I0 (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__I0 (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__I0 (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10737__I (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__I (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__I (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__I (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__I (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__I (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__I (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08321__I (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__I0 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08425__I0 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__I0 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__I0 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__S (.I(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__S (.I(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08328__S (.I(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__S (.I(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__I (.I(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__I (.I(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10411__I (.I(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08326__I (.I(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__I (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__I (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__I (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__I (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__I0 (.I(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08427__I0 (.I(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__I0 (.I(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08328__I0 (.I(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__I (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__I (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__I (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__I (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__I (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__I (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__I (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__I (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__I0 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__I0 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__I0 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__I0 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__I (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__I (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__I (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08337__I (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08471__I0 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__I0 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__I0 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__I0 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__I (.I(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__I (.I(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__I (.I(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__I (.I(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__I (.I(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__I (.I(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08522__I (.I(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08342__I (.I(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__I0 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__I0 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__I0 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__I0 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__S (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__S (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__S (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__S (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__I (.I(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__I (.I(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__I (.I(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__I (.I(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__I (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__I (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__I (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__I (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__I0 (.I(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__I0 (.I(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__I0 (.I(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__I0 (.I(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__I (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__I (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__I (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__I (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__I (.I(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__I (.I(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__I (.I(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__I (.I(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__I0 (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__I0 (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__I0 (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__I0 (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__I (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08702__I (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__I (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__I (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__I0 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__I0 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__I0 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__I0 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__A2 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__A2 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A2 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__I (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__I (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__I (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__I (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__S (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__S (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__S (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__S (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__S (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__S (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__S (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__S (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__S (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__S (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__S (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__S (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__A2 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08433__I (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__I (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__I (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__I (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__S (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__S (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__S (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__S (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08572__A4 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__A3 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__A3 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__A3 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__I (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__I (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__I (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__I (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08453__S (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08451__S (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__S (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08447__S (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__S (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__S (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__S (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__S (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08471__S (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__S (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__S (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__S (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__S (.I(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__S (.I(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__S (.I(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__S (.I(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__I0 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__I0 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__I0 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__I0 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__I (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__I (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__I (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__I (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__S (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__S (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__S (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__S (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__I0 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__I0 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__I0 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__I0 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__I0 (.I(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__I0 (.I(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__I0 (.I(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__I0 (.I(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__I0 (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08580__I0 (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__I0 (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__I0 (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__I0 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08583__I0 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__I0 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__I0 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__I0 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__I0 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__I0 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__I0 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__I0 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__I0 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__I0 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__I0 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__I0 (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__I0 (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__I0 (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__I0 (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__I0 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__I0 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__I0 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__I0 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__S (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__S (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__S (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__S (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__I0 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__I0 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__I0 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__I0 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__I0 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__I0 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__I0 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__I0 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08637__I0 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__I0 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__I0 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__I0 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__I0 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__I0 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__I0 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__I0 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08642__I0 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08603__I0 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__I0 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__I0 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__I0 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08605__I0 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__I0 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__I0 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__I0 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__I0 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__I0 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08533__I0 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__I (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__I (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__I (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__I (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__S (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__S (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__S (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__S (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__S (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__S (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__S (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__S (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__I (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__I (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08582__I (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08573__I (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08580__S (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__S (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__S (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__S (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__S (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__S (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__S (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__S (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__S (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08605__S (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08603__S (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__S (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09321__A3 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__A4 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__A3 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__A3 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__I (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__I (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08621__I (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__I (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__S (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__S (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__S (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__S (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__S (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__S (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__S (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__S (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08637__S (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__S (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__S (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__S (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__I0 (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__I0 (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__I0 (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__I0 (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09188__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08651__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__A1 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__A1 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__A1 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A2 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__I (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__I (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__I (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__I (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__S (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__S (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__S (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__S (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__I0 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__I0 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__I0 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__I0 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__I0 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__I0 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__I0 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__I0 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__I0 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__I0 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__I0 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__I0 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__I0 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__I0 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__I0 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__I0 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__S (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__S (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__S (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__S (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__I0 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__I0 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__I0 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__I0 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__I0 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__I0 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__I0 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__I0 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__I0 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__I0 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__I0 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__I0 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__I0 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__I0 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__I0 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__I0 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__S (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__S (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__S (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__S (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__I0 (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__I0 (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__I0 (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__I0 (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__I0 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__I0 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__I0 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__I0 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__I0 (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__I0 (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08731__I0 (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__I0 (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__I0 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__I0 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__I0 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__I0 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__S (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__S (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08697__S (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__S (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__I0 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__I0 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__I0 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08697__I0 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__I0 (.I(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__I0 (.I(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08738__I0 (.I(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__I0 (.I(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__I0 (.I(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__I0 (.I(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__I0 (.I(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__I0 (.I(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08733__I (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08724__I (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__I (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08706__I (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__S (.I(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__S (.I(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__S (.I(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__S (.I(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__S (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__S (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__S (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__S (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__I (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__I (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__I (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__I (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__S (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__S (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__S (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__S (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__S (.I(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__S (.I(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__S (.I(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__S (.I(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__S (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__S (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__S (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__S (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__S (.I(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__S (.I(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__S (.I(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__S (.I(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__A1 (.I(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A1 (.I(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A1 (.I(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A1 (.I(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09190__I (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__I (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__I (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__I (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__I (.I(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__I (.I(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__I (.I(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__I (.I(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__S (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__S (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__S (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__S (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__S (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__S (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__S (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__S (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__S (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__S (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__S (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__S (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__I0 (.I(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__I0 (.I(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__I0 (.I(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__I0 (.I(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11913__A1 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__A1 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A1 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A2 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08866__I (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__I (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__I (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__I (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__S (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__S (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__S (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__S (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__I0 (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__I0 (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__I0 (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__I0 (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__I0 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__I0 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__I0 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__I0 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__I0 (.I(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__I0 (.I(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__I0 (.I(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__I0 (.I(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__I0 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__I0 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__I0 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__I0 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__S (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__S (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__S (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__S (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__I0 (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__I0 (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__I0 (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__I0 (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__I0 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__I0 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__I0 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__I0 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__I0 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__I0 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08895__I0 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__I0 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__I0 (.I(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08937__I0 (.I(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__I0 (.I(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__I0 (.I(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__S (.I(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__S (.I(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__S (.I(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__S (.I(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__I0 (.I(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__I0 (.I(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__I0 (.I(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__I0 (.I(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__I0 (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__I0 (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__I0 (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__I0 (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__I0 (.I(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__I0 (.I(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__I0 (.I(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__I0 (.I(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__I0 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__I0 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__I0 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__I0 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__S (.I(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__S (.I(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__S (.I(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__S (.I(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__I0 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__I0 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__I0 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__I0 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__I0 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__I0 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__I0 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__I0 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__I0 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__I0 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__I0 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__I0 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__I (.I(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__I (.I(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__I (.I(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__I (.I(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__S (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__S (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__S (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__S (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__S (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__S (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__S (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__S (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__S (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__S (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__S (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__S (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11670__A1 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__A1 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__A1 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__I (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__A1 (.I(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__A1 (.I(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__A1 (.I(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__A1 (.I(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__I (.I(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__I (.I(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__I (.I(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__I (.I(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__S (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__S (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__S (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__S (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__S (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__S (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__S (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08937__S (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__S (.I(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__S (.I(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__S (.I(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__S (.I(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11685__A1 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__A1 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11167__A1 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__I (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10906__A1 (.I(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A1 (.I(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A1 (.I(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__A1 (.I(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__I (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__I (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08966__I (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__I (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__S (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__S (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__S (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__S (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__S (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__S (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__S (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__S (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__I (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__I (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__I (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08994__I (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__I (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__I (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__I (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08995__I (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__I0 (.I(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__I0 (.I(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__I0 (.I(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__I0 (.I(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11699__A1 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11440__A1 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__A1 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__I (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__A1 (.I(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__A1 (.I(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A1 (.I(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A1 (.I(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__I (.I(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__I (.I(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__I (.I(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__I (.I(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__S (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__S (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__S (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__S (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__I (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__I (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__I (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__I (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__I (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09365__I (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09195__I (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__I (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__I0 (.I(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__I0 (.I(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09077__I0 (.I(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__I0 (.I(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__I (.I(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__I (.I(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__I (.I(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__I (.I(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__I (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09368__I (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09198__I (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__I (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__I0 (.I(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__I0 (.I(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__I0 (.I(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__I0 (.I(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__I (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__I (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__I (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__I (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__I (.I(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__I (.I(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__I (.I(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__I (.I(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__I0 (.I(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__I0 (.I(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__I0 (.I(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__I0 (.I(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__I (.I(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__I (.I(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__I (.I(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__I (.I(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__I (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__I (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__I (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__I (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__I0 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09121__I0 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09084__I0 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__I0 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10956__I (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__I (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__I (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__I (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__I (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__I (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__I (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__I (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__I0 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__I0 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09086__I0 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__I0 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__I (.I(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__I (.I(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09211__I (.I(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__I (.I(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__I0 (.I(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__I0 (.I(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09088__I0 (.I(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__I0 (.I(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__I (.I(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09384__I (.I(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__I (.I(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__I (.I(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__I0 (.I(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__I0 (.I(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__I0 (.I(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__I0 (.I(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__I (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__I (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09217__I (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__I (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__I0 (.I(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__I0 (.I(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__I0 (.I(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__I0 (.I(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__S (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__S (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__S (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__S (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__I (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__I (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09221__I (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__I (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__I0 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__I0 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09095__I0 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__I0 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__I (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09394__I (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09224__I (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__I (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__I0 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__I0 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__I0 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__I0 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__I (.I(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__I (.I(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__I (.I(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__I (.I(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__I0 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__I0 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__I0 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__I0 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__I (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__I (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__I (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__I (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09178__I0 (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__I0 (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__I0 (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__I0 (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__I (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__I (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09234__I (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__I (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09180__I0 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__I0 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__I0 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__I0 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09578__I (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__I (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09237__I (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__I (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__I0 (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__I0 (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__I0 (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__I0 (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__I (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__I (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09240__I (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__I (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09184__I0 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__I0 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__I0 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__I0 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11714__A1 (.I(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__A1 (.I(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11197__A1 (.I(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__I (.I(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__A1 (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__A1 (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__A1 (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__A1 (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__I (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__I (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09083__I (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__I (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__S (.I(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__S (.I(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09077__S (.I(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__S (.I(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__S (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__S (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09095__S (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__S (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__S (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__S (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__S (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__S (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__I (.I(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__I (.I(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__I (.I(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__I (.I(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__S (.I(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__S (.I(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__S (.I(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__S (.I(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__S (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__S (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__S (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__S (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__S (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__S (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__S (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__S (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11748__A1 (.I(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11495__A1 (.I(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__A1 (.I(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__I (.I(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__A1 (.I(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__A1 (.I(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09840__A1 (.I(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09149__A1 (.I(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__I (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__I (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__I (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__I (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__S (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__S (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__S (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__S (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__S (.I(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__S (.I(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__S (.I(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__S (.I(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__I0 (.I(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__I0 (.I(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__I0 (.I(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__I0 (.I(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11762__A1 (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11509__A1 (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__A1 (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__I (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10990__A1 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10546__A1 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__A1 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__A1 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__A2 (.I(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09284__A2 (.I(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09245__A2 (.I(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__A2 (.I(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__I (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09218__I (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__I (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__I (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09202__S (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__S (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__S (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__S (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__I0 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__I0 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__I0 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__I0 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__I0 (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09290__I0 (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09251__I0 (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__I0 (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__I0 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__I0 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__I0 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09202__I0 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09334__I0 (.I(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__I0 (.I(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__I0 (.I(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09206__I0 (.I(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__S (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09212__S (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09209__S (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09206__S (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__I0 (.I(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__I0 (.I(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__I0 (.I(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09209__I0 (.I(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09338__I0 (.I(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__I0 (.I(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09260__I0 (.I(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09212__I0 (.I(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09340__I0 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09301__I0 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__I0 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__I0 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__I0 (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__I0 (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09265__I0 (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09219__I0 (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__S (.I(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__S (.I(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__S (.I(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09219__S (.I(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__I0 (.I(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__I0 (.I(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09267__I0 (.I(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__I0 (.I(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__I0 (.I(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__I0 (.I(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09269__I0 (.I(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__I0 (.I(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__I0 (.I(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__I0 (.I(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09271__I0 (.I(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__I0 (.I(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__I0 (.I(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09313__I0 (.I(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09274__I0 (.I(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__I0 (.I(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__I0 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__I0 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__I0 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09235__I0 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__I0 (.I(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__I0 (.I(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09278__I0 (.I(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__I0 (.I(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09358__I0 (.I(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__I0 (.I(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__I0 (.I(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09241__I0 (.I(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11777__A1 (.I(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11524__A1 (.I(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__A1 (.I(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__I (.I(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10598__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09245__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09273__I (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__I (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__I (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__I (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__S (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09251__S (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__S (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__S (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__S (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09260__S (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__S (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__S (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09271__S (.I(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09269__S (.I(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09267__S (.I(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09265__S (.I(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__S (.I(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09278__S (.I(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__S (.I(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09274__S (.I(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11796__A1 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11543__A1 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11284__A1 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09283__I (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__A1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__A1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__A1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09284__A1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09312__I (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__I (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__I (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09285__I (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__S (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09290__S (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__S (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__S (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11811__A1 (.I(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11558__A1 (.I(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__A1 (.I(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09322__I (.I(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11039__A1 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__A1 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10005__A1 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__I (.I(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__I (.I(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__I (.I(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__I (.I(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__S (.I(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__S (.I(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__S (.I(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__S (.I(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__S (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__S (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__S (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__S (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__I0 (.I(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__I0 (.I(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__I0 (.I(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__I0 (.I(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__I (.I(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__I (.I(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09375__I (.I(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__I (.I(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09372__S (.I(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__S (.I(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__S (.I(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__S (.I(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__I0 (.I(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__I0 (.I(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__I0 (.I(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__I0 (.I(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09500__I0 (.I(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__I0 (.I(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__I0 (.I(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__I0 (.I(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__I0 (.I(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__I0 (.I(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__I0 (.I(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09372__I0 (.I(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__I0 (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__I0 (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__I0 (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09376__I0 (.I(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__I0 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__I0 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__I0 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__I0 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__I0 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__I0 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__I0 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09382__I0 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__I0 (.I(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__I0 (.I(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__I0 (.I(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09385__I0 (.I(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__I0 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__I0 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__I0 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__I0 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__S (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__S (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09392__S (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__S (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__I0 (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__I0 (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__I0 (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09392__I0 (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__I0 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__I0 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09439__I0 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__I0 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__I0 (.I(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__I0 (.I(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__I0 (.I(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__I0 (.I(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__I0 (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09483__I0 (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__I0 (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__I0 (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__I0 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__I0 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09446__I0 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__I0 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__I0 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__I0 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__I0 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09408__I0 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__I0 (.I(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09489__I0 (.I(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__I0 (.I(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__I0 (.I(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11840__A1 (.I(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11587__A1 (.I(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11328__A1 (.I(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__I (.I(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11069__A1 (.I(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__A1 (.I(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__A1 (.I(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__A1 (.I(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__I (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__I (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__I (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__I (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__S (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__S (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__S (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__S (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__S (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09439__S (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__S (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__S (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11859__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__I (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__A1 (.I(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11088__A1 (.I(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__A1 (.I(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__A1 (.I(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__I (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09473__I (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__I (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__I (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__S (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__S (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__S (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__S (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__I (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__I (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__I (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__I (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__A2 (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A2 (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A2 (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A2 (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09522__I (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__I (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__I (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__I (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__S (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__S (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__S (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__S (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__S (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__S (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__S (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__S (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__I0 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__I0 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09586__I0 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__I0 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__I (.I(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__I (.I(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__I (.I(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__I (.I(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__S (.I(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__S (.I(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__S (.I(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__S (.I(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__I0 (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__I0 (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__I0 (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__I0 (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__I0 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09627__I0 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__I0 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__I0 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__I0 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__I0 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__I0 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__I0 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__I0 (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__I0 (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__I0 (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__I0 (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__S (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__S (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__S (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__S (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__I0 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__I0 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__I0 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__I0 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__I0 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__I0 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__I0 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__I0 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__I0 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__I0 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__I0 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__I0 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__I0 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__I0 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__I0 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__I0 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__S (.I(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__S (.I(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__S (.I(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__S (.I(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__I0 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__I0 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__I0 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__I0 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__I0 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__I0 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__I0 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__I0 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__I0 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__I0 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__I0 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__I0 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__I0 (.I(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__I0 (.I(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__I0 (.I(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__I0 (.I(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__I0 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__I0 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__I0 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09576__I0 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__I0 (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__I0 (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__I0 (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__I0 (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__I0 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__I0 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09619__I0 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09582__I0 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__I (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__I (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__I (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__I (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__S (.I(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__S (.I(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__S (.I(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09586__S (.I(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__S (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__S (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__S (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__S (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__S (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__S (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__S (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__S (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__I (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__I (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__I (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__I (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__S (.I(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09627__S (.I(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__S (.I(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__S (.I(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__S (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__S (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__S (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__S (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__S (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__S (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__S (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__S (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__I (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__I (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09669__I (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__I (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__S (.I(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__S (.I(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__S (.I(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__S (.I(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__S (.I(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__S (.I(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__S (.I(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__S (.I(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__S (.I(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__S (.I(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__S (.I(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__S (.I(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__I0 (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__I0 (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__I0 (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__I0 (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__I (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__I (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__I (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__I (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__S (.I(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__S (.I(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__S (.I(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__S (.I(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__I0 (.I(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__I0 (.I(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__I0 (.I(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__I0 (.I(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__I0 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__I0 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__I0 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__I0 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__I0 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__I0 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__I0 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__I0 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__I0 (.I(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__I0 (.I(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09776__I0 (.I(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__I0 (.I(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10227__I (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__I (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__I (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__I (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__I0 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__I0 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__I0 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__I0 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__I0 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__I0 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__I0 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__I0 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__I (.I(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__I (.I(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__I (.I(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09728__I (.I(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__I0 (.I(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__I0 (.I(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__I0 (.I(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__I0 (.I(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__I0 (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__I0 (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__I0 (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__I0 (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__S (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__S (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__S (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__S (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__I0 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__I0 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__I0 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__I0 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09864__I0 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__I0 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__I0 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__I0 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__I0 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09828__I0 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__I0 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__I0 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__I0 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__I0 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__I0 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__I0 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__I0 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__I0 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09796__I0 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09755__I0 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__I0 (.I(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__I0 (.I(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__I0 (.I(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__I0 (.I(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__I0 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__I0 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__I0 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__I0 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09793__I (.I(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__I (.I(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__I (.I(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09766__I (.I(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__S (.I(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__S (.I(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__S (.I(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__S (.I(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__S (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__S (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__S (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__S (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__S (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__S (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09796__S (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__S (.I(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__I (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09821__I (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__I (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__I (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__S (.I(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__S (.I(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__S (.I(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__S (.I(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09828__S (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__S (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__S (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__S (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__S (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__S (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__S (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__S (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__A2 (.I(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__A2 (.I(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__A2 (.I(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09840__A2 (.I(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__I (.I(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__I (.I(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09850__I (.I(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__I (.I(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__S (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__S (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__S (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__S (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__S (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__S (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__S (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__S (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__S (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09864__S (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__S (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__S (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__I0 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__I0 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__I0 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__I0 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__I (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__I (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__I (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__I (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__S (.I(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09886__S (.I(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__S (.I(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__S (.I(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__I0 (.I(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__I0 (.I(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__I0 (.I(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__I0 (.I(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__I0 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__I0 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__I0 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09886__I0 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__I0 (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__I0 (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__I0 (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__I0 (.I(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__I0 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__I0 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09941__I0 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__I0 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__I0 (.I(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09980__I0 (.I(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__I0 (.I(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__I0 (.I(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__I0 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__I0 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__I0 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__I0 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__I0 (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__I0 (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09947__I0 (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09902__I0 (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__I0 (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__I0 (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__I0 (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__I0 (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__I0 (.I(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__I0 (.I(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__I0 (.I(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__I0 (.I(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__I0 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__I0 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__I0 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__I0 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__I0 (.I(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09993__I0 (.I(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__I0 (.I(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__I0 (.I(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__I0 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__I0 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09959__I0 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__I0 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__I0 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__I0 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__I0 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__I0 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__I0 (.I(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__I0 (.I(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09963__I0 (.I(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__I0 (.I(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__I0 (.I(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__I0 (.I(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__I0 (.I(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__I0 (.I(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__I (.I(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__I (.I(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__I (.I(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__I (.I(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__S (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__S (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__S (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__S (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__S (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__S (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__S (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__S (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__S (.I(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09963__S (.I(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__S (.I(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09959__S (.I(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__I (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__I (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__I (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__I (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__S (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__S (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__S (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__S (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09993__S (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__S (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__S (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__S (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__S (.I(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__S (.I(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__S (.I(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__S (.I(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__A2 (.I(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__A2 (.I(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__A2 (.I(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10005__A2 (.I(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__I (.I(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10024__I (.I(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10015__I (.I(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__I (.I(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__S (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__S (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__S (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__S (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__S (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__S (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__S (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__S (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__S (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__S (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__S (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__S (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__S (.I(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__S (.I(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__S (.I(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__S (.I(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__I0 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__I0 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__I0 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10045__I0 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__I (.I(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__I (.I(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__I (.I(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__I (.I(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__S (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__S (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__S (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10045__S (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__I0 (.I(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__I0 (.I(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__I0 (.I(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__I0 (.I(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__I0 (.I(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__I0 (.I(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__I0 (.I(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__I0 (.I(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__I0 (.I(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10140__I0 (.I(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__I0 (.I(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__I0 (.I(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__I0 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__I0 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__I0 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__I0 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__I0 (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__I0 (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__I0 (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__I0 (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__I0 (.I(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__I0 (.I(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__I0 (.I(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__I0 (.I(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__I0 (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__I0 (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__I0 (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__I0 (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__I0 (.I(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__I0 (.I(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__I0 (.I(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__I0 (.I(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__S (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__S (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__S (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__S (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__I0 (.I(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__I0 (.I(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__I0 (.I(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__I0 (.I(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__I0 (.I(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__I0 (.I(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__I0 (.I(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__I0 (.I(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__I0 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__I0 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__I0 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__I0 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__I0 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10161__I0 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__I0 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__I0 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__I0 (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__I0 (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__I0 (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__I0 (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__I0 (.I(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__I0 (.I(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__I0 (.I(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__I0 (.I(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__I0 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__I0 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__I0 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__I0 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__I (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__I (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__I (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__I (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__S (.I(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__S (.I(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__S (.I(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__S (.I(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__S (.I(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__S (.I(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__S (.I(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__S (.I(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__S (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__S (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__S (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__S (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__S (.I(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__S (.I(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__S (.I(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__S (.I(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__I (.I(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__I (.I(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__I (.I(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10133__I (.I(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10140__S (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__S (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__S (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__S (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__S (.I(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__S (.I(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__S (.I(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__S (.I(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__S (.I(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__S (.I(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__S (.I(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10161__S (.I(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10672__I (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__I (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__I (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__I (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__A2 (.I(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__A2 (.I(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__A2 (.I(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A2 (.I(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__I (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__I (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__I (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__I (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__S (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__S (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__S (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__S (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__S (.I(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__S (.I(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__S (.I(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__S (.I(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__S (.I(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__S (.I(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__S (.I(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__S (.I(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__I0 (.I(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__I0 (.I(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__I0 (.I(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__I0 (.I(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__I (.I(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__I (.I(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__I (.I(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10211__I (.I(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__S (.I(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__S (.I(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__S (.I(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__S (.I(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__I0 (.I(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__I0 (.I(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__I0 (.I(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__I0 (.I(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__I0 (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__I0 (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__I0 (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__I0 (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__I0 (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__I0 (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__I0 (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__I0 (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__I0 (.I(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__I0 (.I(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__I0 (.I(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__I0 (.I(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__S (.I(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__S (.I(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__S (.I(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__S (.I(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__I0 (.I(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__I0 (.I(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__I0 (.I(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__I0 (.I(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__I0 (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__I0 (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__I0 (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__I0 (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__I0 (.I(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__I0 (.I(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__I0 (.I(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__I0 (.I(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10357__I0 (.I(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__I0 (.I(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__I0 (.I(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__I0 (.I(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__S (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__S (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__S (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__S (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__I0 (.I(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__I0 (.I(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__I0 (.I(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__I0 (.I(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__I0 (.I(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__I0 (.I(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__I0 (.I(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__I0 (.I(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__I0 (.I(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__I0 (.I(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__I0 (.I(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__I0 (.I(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__I0 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__I0 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__I0 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__I0 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__I0 (.I(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__I0 (.I(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__I0 (.I(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__I0 (.I(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__I0 (.I(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__I0 (.I(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__I0 (.I(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__I0 (.I(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__I0 (.I(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__I0 (.I(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__I0 (.I(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__I0 (.I(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__I (.I(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__I (.I(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__I (.I(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__I (.I(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__S (.I(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__S (.I(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__S (.I(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__S (.I(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__S (.I(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__S (.I(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__S (.I(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__S (.I(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__S (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__S (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__S (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__S (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__I (.I(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__I (.I(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10309__I (.I(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__I (.I(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__S (.I(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__S (.I(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__S (.I(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__S (.I(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__S (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__S (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__S (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__S (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__S (.I(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__S (.I(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__S (.I(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__S (.I(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__S (.I(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__S (.I(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__S (.I(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__S (.I(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__A2 (.I(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__A2 (.I(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__A2 (.I(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A2 (.I(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__I (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__I (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__I (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__I (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__S (.I(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__S (.I(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__S (.I(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__S (.I(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__S (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__S (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__S (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10357__S (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__I (.I(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10710__I (.I(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__I (.I(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__I (.I(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__I0 (.I(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10472__I0 (.I(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__I0 (.I(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__I0 (.I(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__I (.I(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__I (.I(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10394__I (.I(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__I (.I(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__S (.I(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__S (.I(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__S (.I(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__S (.I(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10876__I (.I(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10715__I (.I(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__I (.I(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__I (.I(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__I0 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10474__I0 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__I0 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__I0 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__I (.I(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__I (.I(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__I (.I(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10385__I (.I(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__I0 (.I(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__I0 (.I(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__I0 (.I(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__I0 (.I(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__I (.I(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__I (.I(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10556__I (.I(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__I (.I(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__I0 (.I(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__I0 (.I(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__I0 (.I(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__I0 (.I(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__I (.I(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__I (.I(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__I (.I(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__I (.I(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__I0 (.I(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10481__I0 (.I(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__I0 (.I(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__I0 (.I(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__S (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__S (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__S (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__S (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__I (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10728__I (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__I (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10398__I (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__I0 (.I(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__I0 (.I(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__I0 (.I(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__I0 (.I(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10523__I0 (.I(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__I0 (.I(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__I0 (.I(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__I0 (.I(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__I0 (.I(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10487__I0 (.I(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__I0 (.I(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__I0 (.I(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__I0 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__I0 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__I0 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__I0 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__S (.I(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10415__S (.I(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10412__S (.I(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__S (.I(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10530__I0 (.I(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__I0 (.I(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__I0 (.I(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10412__I0 (.I(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__I0 (.I(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__I0 (.I(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__I0 (.I(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10415__I0 (.I(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10534__I0 (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__I0 (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__I0 (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__I0 (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10537__I0 (.I(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__I0 (.I(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10462__I0 (.I(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10422__I0 (.I(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10539__I0 (.I(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10501__I0 (.I(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__I0 (.I(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__I0 (.I(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10541__I0 (.I(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__I0 (.I(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__I0 (.I(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10428__I0 (.I(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__I0 (.I(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__I0 (.I(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__I0 (.I(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__I0 (.I(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__I (.I(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__I (.I(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__I (.I(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__I (.I(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__S (.I(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__S (.I(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__S (.I(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__S (.I(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__S (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__S (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__S (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__S (.I(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__S (.I(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__S (.I(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__S (.I(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__S (.I(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__S (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__S (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__S (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10462__S (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10498__I (.I(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__I (.I(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__I (.I(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10471__I (.I(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__S (.I(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__S (.I(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10474__S (.I(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10472__S (.I(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10487__S (.I(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__S (.I(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__S (.I(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10481__S (.I(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__S (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__S (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__S (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__S (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__S (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__S (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10501__S (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__S (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10536__I (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__I (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__I (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10509__I (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__S (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__S (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__S (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__S (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__S (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10523__S (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__S (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__S (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10534__S (.I(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__S (.I(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10530__S (.I(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__S (.I(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10675__I0 (.I(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10637__I0 (.I(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__I0 (.I(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__I0 (.I(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10586__I (.I(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__I (.I(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__I (.I(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__I (.I(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__S (.I(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10554__S (.I(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__S (.I(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__S (.I(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__I0 (.I(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10639__I0 (.I(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__I0 (.I(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__I0 (.I(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__I0 (.I(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__I0 (.I(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__I0 (.I(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10554__I0 (.I(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10681__I0 (.I(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__I0 (.I(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10606__I0 (.I(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__I0 (.I(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10684__I0 (.I(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__I0 (.I(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10609__I0 (.I(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__I0 (.I(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__I0 (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10648__I0 (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__I0 (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10564__I0 (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10688__I0 (.I(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__I0 (.I(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__I0 (.I(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10567__I0 (.I(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__I0 (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__I0 (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__I0 (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__I0 (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10693__I0 (.I(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__I0 (.I(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10618__I0 (.I(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__I0 (.I(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__S (.I(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__S (.I(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__S (.I(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__S (.I(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__I0 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__I0 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10620__I0 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__I0 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__I0 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__I0 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__I0 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__I0 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10699__I0 (.I(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10661__I0 (.I(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__I0 (.I(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__I0 (.I(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10702__I0 (.I(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__I0 (.I(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__I0 (.I(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__I0 (.I(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__I0 (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__I0 (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10629__I0 (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10590__I0 (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10706__I0 (.I(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10668__I0 (.I(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10631__I0 (.I(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__I0 (.I(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__I0 (.I(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__I0 (.I(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__I0 (.I(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__I0 (.I(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__I (.I(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10617__I (.I(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10608__I (.I(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10599__I (.I(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10606__S (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__S (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__S (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__S (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__S (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__S (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10620__S (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10618__S (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__I (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10654__I (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__I (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__I (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__S (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__S (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10639__S (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10637__S (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__S (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__S (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10648__S (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__S (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10661__S (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__S (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__S (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__S (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10701__I (.I(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10692__I (.I(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10683__I (.I(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10674__I (.I(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10681__S (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__S (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__S (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10675__S (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__S (.I(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10688__S (.I(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__S (.I(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10684__S (.I(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10699__S (.I(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__S (.I(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__S (.I(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10693__S (.I(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__I0 (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__I0 (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10765__I0 (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__I0 (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__I (.I(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10738__I (.I(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10725__I (.I(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__I (.I(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__S (.I(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__S (.I(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__S (.I(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__S (.I(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__I0 (.I(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__I0 (.I(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__I0 (.I(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__I0 (.I(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__I0 (.I(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10847__I0 (.I(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__I0 (.I(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__I0 (.I(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__I0 (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10849__I0 (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__I0 (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__I0 (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__I0 (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__I0 (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__I0 (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__I0 (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__S (.I(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10732__S (.I(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10729__S (.I(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__S (.I(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10868__I0 (.I(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10853__I0 (.I(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__I0 (.I(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10729__I0 (.I(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11967__I0 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11928__I0 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__I0 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10732__I0 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11969__I0 (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11930__I0 (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__I0 (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__I0 (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11971__I0 (.I(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11933__I0 (.I(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__I0 (.I(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__I0 (.I(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__S (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__S (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__S (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__S (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11973__I0 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11935__I0 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__I0 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__I0 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11976__I0 (.I(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11937__I0 (.I(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10787__I0 (.I(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__I0 (.I(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11978__I0 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11939__I0 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__I0 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__I0 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11980__I0 (.I(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11942__I0 (.I(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10792__I0 (.I(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__I0 (.I(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11982__I0 (.I(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11944__I0 (.I(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10794__I0 (.I(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__I0 (.I(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11984__I0 (.I(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11946__I0 (.I(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__I0 (.I(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__I0 (.I(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11948__I0 (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10835__I1 (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__I0 (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__I0 (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__I (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__I (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10773__I (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__I (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__S (.I(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__S (.I(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__S (.I(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10765__S (.I(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__S (.I(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__S (.I(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__S (.I(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__S (.I(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__S (.I(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10787__S (.I(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__S (.I(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__S (.I(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10828__I (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10819__I (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__I (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__I (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__S (.I(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__S (.I(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__S (.I(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__S (.I(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__S (.I(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10824__S (.I(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__S (.I(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10820__S (.I(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11038__I (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__I (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__I (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10840__I (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10853__S (.I(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__S (.I(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10842__I (.I(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10849__S (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10847__S (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__S (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__S (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11636__A1 (.I(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11377__A1 (.I(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__A1 (.I(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__A1 (.I(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10868__S (.I(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__S (.I(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10857__I (.I(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__S (.I(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__S (.I(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__S (.I(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__S (.I(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__I0 (.I(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__I0 (.I(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__I0 (.I(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10874__I0 (.I(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11651__A1 (.I(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11392__A1 (.I(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11133__A1 (.I(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__A1 (.I(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__S (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10886__S (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__I (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__S (.I(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10880__S (.I(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__S (.I(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10874__S (.I(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__I0 (.I(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__I0 (.I(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__I0 (.I(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__I0 (.I(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__I0 (.I(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__I0 (.I(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__I0 (.I(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10880__I0 (.I(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__I0 (.I(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__I0 (.I(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__I0 (.I(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10886__I0 (.I(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__I0 (.I(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__I0 (.I(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__I0 (.I(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__I0 (.I(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__S (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__S (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__I (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__S (.I(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__S (.I(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__S (.I(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__S (.I(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__S (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__S (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__I (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__S (.I(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__S (.I(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__S (.I(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__S (.I(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__S (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__S (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__I (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__S (.I(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__S (.I(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__S (.I(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__S (.I(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__I (.I(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11068__I (.I(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11004__I (.I(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__I (.I(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__I0 (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__I0 (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10963__I0 (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__I0 (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__S (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__S (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__I (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__S (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__S (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__S (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__S (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11137__I (.I(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11073__I (.I(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__I (.I(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__I (.I(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__I0 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__I0 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__I0 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__I0 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11140__I (.I(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__I (.I(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__I (.I(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__I (.I(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__I0 (.I(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__I0 (.I(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__I0 (.I(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__I0 (.I(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11143__I (.I(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11079__I (.I(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__I (.I(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__I (.I(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__I0 (.I(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__I0 (.I(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__I0 (.I(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__I0 (.I(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11146__I (.I(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__I (.I(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__I (.I(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__I (.I(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__I0 (.I(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10986__I0 (.I(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__I0 (.I(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__I0 (.I(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11149__I (.I(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11085__I (.I(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__I (.I(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10957__I (.I(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11733__A1 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11480__A1 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__A1 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__A1 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__S (.I(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__S (.I(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__I (.I(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__S (.I(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__S (.I(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__S (.I(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10963__S (.I(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__S (.I(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10986__S (.I(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__I (.I(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__S (.I(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__S (.I(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__S (.I(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__S (.I(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__S (.I(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__S (.I(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10991__I (.I(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__S (.I(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__S (.I(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__S (.I(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__S (.I(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__I0 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11041__I0 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__I0 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__I0 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11022__S (.I(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11019__S (.I(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__I (.I(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__S (.I(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__S (.I(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__S (.I(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__S (.I(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11058__I0 (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__I0 (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__I0 (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__I0 (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__I0 (.I(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__I0 (.I(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__I0 (.I(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__I0 (.I(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11062__I0 (.I(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__I0 (.I(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__I0 (.I(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__I0 (.I(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__I0 (.I(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__I0 (.I(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__I0 (.I(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11022__I0 (.I(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__S (.I(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11034__S (.I(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__I (.I(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__S (.I(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__S (.I(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__S (.I(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__S (.I(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__S (.I(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__S (.I(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__I (.I(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__S (.I(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__S (.I(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__S (.I(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11041__S (.I(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11825__A1 (.I(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__A1 (.I(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__A1 (.I(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__A1 (.I(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__S (.I(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__S (.I(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11055__I (.I(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11062__S (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__S (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11058__S (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__S (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__I0 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__I0 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11090__I0 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__I0 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11086__S (.I(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__S (.I(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11070__I (.I(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__S (.I(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11077__S (.I(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__S (.I(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__S (.I(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11122__I0 (.I(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__I0 (.I(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__I0 (.I(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__I0 (.I(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11124__I0 (.I(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11110__I0 (.I(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__I0 (.I(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11077__I0 (.I(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__I0 (.I(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__I0 (.I(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11096__I0 (.I(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__I0 (.I(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11128__I0 (.I(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__I0 (.I(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__I0 (.I(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__I0 (.I(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__I0 (.I(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__I0 (.I(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11100__I0 (.I(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11086__I0 (.I(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11100__S (.I(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__S (.I(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__I (.I(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11096__S (.I(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__S (.I(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__S (.I(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11090__S (.I(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11298__I (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11235__I (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11166__I (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11103__I (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__A2 (.I(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11133__A2 (.I(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__A2 (.I(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11104__A2 (.I(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__S (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11110__S (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__S (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__S (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__S (.I(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11124__S (.I(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11122__S (.I(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__S (.I(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11183__I0 (.I(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__I0 (.I(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11154__I0 (.I(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11135__I0 (.I(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__S (.I(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__S (.I(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11134__I (.I(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__S (.I(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__S (.I(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__S (.I(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11135__S (.I(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__I0 (.I(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__I0 (.I(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11156__I0 (.I(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__I0 (.I(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__I0 (.I(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__I0 (.I(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__I0 (.I(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__I0 (.I(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11189__I0 (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__I0 (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11160__I0 (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__I0 (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__I0 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__I0 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__I0 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__I0 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11193__I0 (.I(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11179__I0 (.I(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__I0 (.I(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__I0 (.I(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__S (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__S (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__I (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__A2 (.I(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11197__A2 (.I(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__A2 (.I(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11167__A2 (.I(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11179__S (.I(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__S (.I(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__I (.I(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__S (.I(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__S (.I(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__S (.I(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__S (.I(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11189__S (.I(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__S (.I(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__S (.I(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11183__S (.I(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11391__I (.I(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__I (.I(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__I (.I(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__I (.I(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__S (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__S (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__I (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__S (.I(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11207__S (.I(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__S (.I(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__S (.I(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__I (.I(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__I (.I(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__I (.I(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__I (.I(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11399__I (.I(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__I (.I(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__I (.I(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11206__I (.I(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11402__I (.I(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__I (.I(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11275__I (.I(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__I (.I(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11405__I (.I(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11341__I (.I(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11278__I (.I(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11214__I (.I(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11260__I0 (.I(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11246__I0 (.I(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11231__I0 (.I(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__I0 (.I(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__I (.I(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__I (.I(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__I (.I(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11218__I (.I(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__I0 (.I(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11248__I0 (.I(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__I0 (.I(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__I0 (.I(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__S (.I(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11231__S (.I(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11222__I (.I(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11229__S (.I(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11227__S (.I(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__S (.I(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11223__S (.I(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11248__S (.I(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11246__S (.I(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__I (.I(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11244__S (.I(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__S (.I(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__S (.I(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11238__S (.I(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__S (.I(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11260__S (.I(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__I (.I(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__S (.I(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__S (.I(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__S (.I(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__S (.I(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11315__I0 (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__I0 (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__I0 (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11267__I0 (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11282__S (.I(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__S (.I(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11266__I (.I(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__S (.I(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__S (.I(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__S (.I(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11267__S (.I(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__I0 (.I(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__I0 (.I(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__I0 (.I(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__I0 (.I(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__I0 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__I0 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__I0 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__I0 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__I0 (.I(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__I0 (.I(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11292__I0 (.I(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__I0 (.I(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11323__I0 (.I(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__I0 (.I(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11294__I0 (.I(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__I0 (.I(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__I0 (.I(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11311__I0 (.I(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__I0 (.I(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11282__I0 (.I(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__S (.I(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11294__S (.I(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__I (.I(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11311__S (.I(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__S (.I(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11300__I (.I(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__S (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__S (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__S (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__S (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__S (.I(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11323__S (.I(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11314__I (.I(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__S (.I(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__S (.I(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__S (.I(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11315__S (.I(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__I0 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11365__I0 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__I0 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11330__I0 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__S (.I(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11342__S (.I(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11329__I (.I(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__S (.I(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__S (.I(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__S (.I(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11330__S (.I(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11381__I0 (.I(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11367__I0 (.I(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11351__I0 (.I(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__I0 (.I(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11383__I0 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__I0 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__I0 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__I0 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__I0 (.I(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11371__I0 (.I(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__I0 (.I(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__I0 (.I(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__I0 (.I(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11373__I0 (.I(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11357__I0 (.I(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11342__I0 (.I(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11389__I0 (.I(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11375__I0 (.I(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__I0 (.I(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__I0 (.I(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__S (.I(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11357__S (.I(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__I (.I(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__S (.I(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__S (.I(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11351__S (.I(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__S (.I(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11557__I (.I(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11494__I (.I(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11425__I (.I(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__I (.I(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__A2 (.I(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11392__A2 (.I(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11377__A2 (.I(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11363__A2 (.I(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11375__S (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11373__S (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11364__I (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11389__S (.I(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__S (.I(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11378__I (.I(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__S (.I(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11383__S (.I(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11381__S (.I(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__S (.I(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__I0 (.I(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11428__I0 (.I(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__I0 (.I(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__I0 (.I(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__S (.I(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11406__S (.I(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11393__I (.I(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__S (.I(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11400__S (.I(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__S (.I(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__S (.I(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11444__I0 (.I(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11430__I0 (.I(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__I0 (.I(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__I0 (.I(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11446__I0 (.I(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11432__I0 (.I(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__I0 (.I(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11400__I0 (.I(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__I0 (.I(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__I0 (.I(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__I0 (.I(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__I0 (.I(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11450__I0 (.I(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11436__I0 (.I(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__I0 (.I(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11406__I0 (.I(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__I0 (.I(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11438__I0 (.I(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11423__I0 (.I(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__I0 (.I(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11423__S (.I(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__S (.I(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__I (.I(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__S (.I(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__S (.I(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__S (.I(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__S (.I(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11480__A2 (.I(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__A2 (.I(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11440__A2 (.I(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__A2 (.I(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11438__S (.I(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11436__S (.I(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11427__I (.I(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__S (.I(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11450__S (.I(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11441__I (.I(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__S (.I(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11446__S (.I(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11444__S (.I(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__S (.I(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11511__I0 (.I(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11497__I0 (.I(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__I0 (.I(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11458__I0 (.I(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11655__I (.I(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11591__I (.I(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11528__I (.I(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11461__I (.I(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11513__I0 (.I(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11499__I0 (.I(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11484__I0 (.I(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11462__I0 (.I(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__I0 (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11501__I0 (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11486__I0 (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__I0 (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11517__I0 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11503__I0 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__I0 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11470__I0 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11664__I (.I(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11600__I (.I(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11537__I (.I(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11473__I (.I(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11519__I0 (.I(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11505__I0 (.I(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11490__I0 (.I(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11474__I0 (.I(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11521__I0 (.I(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11507__I0 (.I(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11492__I0 (.I(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11478__I0 (.I(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11492__S (.I(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11490__S (.I(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11481__I (.I(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__S (.I(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11486__S (.I(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11484__S (.I(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__S (.I(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11543__A2 (.I(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11524__A2 (.I(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11509__A2 (.I(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11495__A2 (.I(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11507__S (.I(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11505__S (.I(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11496__I (.I(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11503__S (.I(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11501__S (.I(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11499__S (.I(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11497__S (.I(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11517__S (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__S (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11513__S (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11511__S (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11574__I0 (.I(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11560__I0 (.I(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11545__I0 (.I(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11526__I0 (.I(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11541__S (.I(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11538__S (.I(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11525__I (.I(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__S (.I(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11532__S (.I(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11529__S (.I(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11526__S (.I(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11576__I0 (.I(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11562__I0 (.I(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11547__I0 (.I(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11529__I0 (.I(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__I0 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11564__I0 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11549__I0 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11532__I0 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__I0 (.I(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11566__I0 (.I(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__I0 (.I(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__I0 (.I(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11582__I0 (.I(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11568__I0 (.I(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11553__I0 (.I(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11538__I0 (.I(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11584__I0 (.I(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11570__I0 (.I(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11555__I0 (.I(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11541__I0 (.I(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__S (.I(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11549__S (.I(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11547__S (.I(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11545__S (.I(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__A2 (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11587__A2 (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__A2 (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11558__A2 (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11570__S (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11568__S (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11559__I (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11566__S (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11564__S (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11562__S (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11560__S (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11584__S (.I(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11582__S (.I(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11573__I (.I(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__S (.I(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__S (.I(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11576__S (.I(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11574__S (.I(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11638__I0 (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11624__I0 (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11608__I0 (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11589__I0 (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11604__S (.I(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11601__S (.I(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11588__I (.I(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11598__S (.I(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11595__S (.I(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11592__S (.I(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11589__S (.I(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__I0 (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__I0 (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11610__I0 (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11592__I0 (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__I0 (.I(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11628__I0 (.I(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11612__I0 (.I(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11595__I0 (.I(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11644__I0 (.I(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11630__I0 (.I(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11614__I0 (.I(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11598__I0 (.I(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11646__I0 (.I(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11632__I0 (.I(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11616__I0 (.I(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11601__I0 (.I(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11648__I0 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11634__I0 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11618__I0 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11604__I0 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11618__S (.I(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11616__S (.I(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11607__I (.I(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11614__S (.I(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11612__S (.I(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11610__S (.I(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11608__S (.I(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11810__I (.I(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11747__I (.I(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11684__I (.I(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11621__I (.I(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11670__A2 (.I(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11651__A2 (.I(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11636__A2 (.I(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11622__A2 (.I(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11634__S (.I(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11632__S (.I(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11623__I (.I(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11630__S (.I(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11628__S (.I(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__S (.I(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11624__S (.I(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11648__S (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11646__S (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11637__I (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11644__S (.I(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__S (.I(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__S (.I(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11638__S (.I(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11701__I0 (.I(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11687__I0 (.I(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11672__I0 (.I(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11653__I0 (.I(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11668__S (.I(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11665__S (.I(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11652__I (.I(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11662__S (.I(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11659__S (.I(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11656__S (.I(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11653__S (.I(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11703__I0 (.I(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11689__I0 (.I(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11674__I0 (.I(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11656__I0 (.I(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11705__I0 (.I(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11691__I0 (.I(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11676__I0 (.I(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11659__I0 (.I(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11707__I0 (.I(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11693__I0 (.I(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11678__I0 (.I(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11662__I0 (.I(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11709__I0 (.I(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11695__I0 (.I(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11680__I0 (.I(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11665__I0 (.I(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11711__I0 (.I(_05798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11697__I0 (.I(_05798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11682__I0 (.I(_05798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11668__I0 (.I(_05798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11682__S (.I(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11680__S (.I(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11671__I (.I(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11678__S (.I(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11676__S (.I(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11674__S (.I(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11672__S (.I(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11733__A2 (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11714__A2 (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11699__A2 (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11685__A2 (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11697__S (.I(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11695__S (.I(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11686__I (.I(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11711__S (.I(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11709__S (.I(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11700__I (.I(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11764__I0 (.I(_05825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11750__I0 (.I(_05825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11735__I0 (.I(_05825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11716__I0 (.I(_05825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11766__I0 (.I(_05829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11752__I0 (.I(_05829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11737__I0 (.I(_05829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11719__I0 (.I(_05829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11768__I0 (.I(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11754__I0 (.I(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11739__I0 (.I(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11722__I0 (.I(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11770__I0 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11756__I0 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11741__I0 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11725__I0 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11772__I0 (.I(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11758__I0 (.I(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11743__I0 (.I(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11728__I0 (.I(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11774__I0 (.I(_05837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11760__I0 (.I(_05837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11745__I0 (.I(_05837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11731__I0 (.I(_05837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11741__S (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11739__S (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11737__S (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11735__S (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11796__A2 (.I(_05847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11777__A2 (.I(_05847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11762__A2 (.I(_05847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11748__A2 (.I(_05847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11760__S (.I(_05848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11758__S (.I(_05848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11749__I (.I(_05848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11756__S (.I(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11754__S (.I(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11752__S (.I(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11750__S (.I(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11770__S (.I(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11768__S (.I(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11766__S (.I(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11764__S (.I(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11827__I0 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11813__I0 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11798__I0 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11779__I0 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11794__S (.I(_05865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11791__S (.I(_05865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11778__I (.I(_05865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11788__S (.I(_05866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11785__S (.I(_05866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11782__S (.I(_05866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11779__S (.I(_05866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11829__I0 (.I(_05868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11815__I0 (.I(_05868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11800__I0 (.I(_05868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11782__I0 (.I(_05868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11831__I0 (.I(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11817__I0 (.I(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11802__I0 (.I(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11785__I0 (.I(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11833__I0 (.I(_05872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11819__I0 (.I(_05872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11804__I0 (.I(_05872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11788__I0 (.I(_05872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11835__I0 (.I(_05874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11821__I0 (.I(_05874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11806__I0 (.I(_05874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11791__I0 (.I(_05874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11837__I0 (.I(_05876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11823__I0 (.I(_05876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11808__I0 (.I(_05876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11794__I0 (.I(_05876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11808__S (.I(_05878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11806__S (.I(_05878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11797__I (.I(_05878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11804__S (.I(_05879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11802__S (.I(_05879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11800__S (.I(_05879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11798__S (.I(_05879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11823__S (.I(_05887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11821__S (.I(_05887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11812__I (.I(_05887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11819__S (.I(_05888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11817__S (.I(_05888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11815__S (.I(_05888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11813__S (.I(_05888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11837__S (.I(_05895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11835__S (.I(_05895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11826__I (.I(_05895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11833__S (.I(_05896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11831__S (.I(_05896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11829__S (.I(_05896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11827__S (.I(_05896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11953__I0 (.I(_05903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11915__I0 (.I(_05903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11861__I0 (.I(_05903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11842__I0 (.I(_05903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11857__S (.I(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11854__S (.I(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11841__I (.I(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11851__S (.I(_05905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11848__S (.I(_05905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11845__S (.I(_05905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11842__S (.I(_05905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11955__I0 (.I(_05907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11917__I0 (.I(_05907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11863__I0 (.I(_05907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11845__I0 (.I(_05907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11958__I0 (.I(_05909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11919__I0 (.I(_05909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11865__I0 (.I(_05909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11848__I0 (.I(_05909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11960__I0 (.I(_05911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11921__I0 (.I(_05911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11867__I0 (.I(_05911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11851__I0 (.I(_05911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11962__I0 (.I(_05913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11924__I0 (.I(_05913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11869__I0 (.I(_05913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11854__I0 (.I(_05913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11964__I0 (.I(_05915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11926__I0 (.I(_05915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11871__I0 (.I(_05915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11857__I0 (.I(_05915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11950__A2 (.I(_05926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11913__A2 (.I(_05926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11875__A2 (.I(_05926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11900__I (.I(_05927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11876__I (.I(_05927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11909__S (.I(_05928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11891__I (.I(_05928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11882__I (.I(_05928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11877__I (.I(_05928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11889__S (.I(_05932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11887__S (.I(_05932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11885__S (.I(_05932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11883__S (.I(_05932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11898__S (.I(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11896__S (.I(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11894__S (.I(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11892__S (.I(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11907__S (.I(_05942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11905__S (.I(_05942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11903__S (.I(_05942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11901__S (.I(_05942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11941__I (.I(_05949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11932__I (.I(_05949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11923__I (.I(_05949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11914__I (.I(_05949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11921__S (.I(_05950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11919__S (.I(_05950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11917__S (.I(_05950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11915__S (.I(_05950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11930__S (.I(_05955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11928__S (.I(_05955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11926__S (.I(_05955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11924__S (.I(_05955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11948__S (.I(_05965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11946__S (.I(_05965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11944__S (.I(_05965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11942__S (.I(_05965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11975__I (.I(_05970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11951__I (.I(_05970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11984__S (.I(_05971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11966__I (.I(_05971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11957__I (.I(_05971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11952__I (.I(_05971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11987__A2 (.I(_05972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11986__A2 (.I(_05972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11955__S (.I(_05972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11953__S (.I(_05972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11964__S (.I(_05975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11962__S (.I(_05975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11960__S (.I(_05975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11958__S (.I(_05975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11973__S (.I(_05980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11971__S (.I(_05980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11969__S (.I(_05980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11967__S (.I(_05980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11982__S (.I(_05985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11980__S (.I(_05985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11978__S (.I(_05985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11976__S (.I(_05985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12110__D (.I(_05992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clock_I (.I(clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clock_a_I (.I(clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(col_select_a[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(col_select_a[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(col_select_a[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(col_select_a[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(col_select_a[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(col_select_a[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06066__I (.I(\col_select_trans[0].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06055__I (.I(\col_select_trans[0].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06039__A1 (.I(\col_select_trans[0].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__I (.I(\col_select_trans[1].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06056__A2 (.I(\col_select_trans[1].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06039__A2 (.I(\col_select_trans[1].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06077__I (.I(\col_select_trans[2].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06051__I (.I(\col_select_trans[2].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06041__A1 (.I(\col_select_trans[2].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06061__I (.I(\col_select_trans[3].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06052__I (.I(\col_select_trans[3].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06041__A2 (.I(\col_select_trans[3].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12046__D (.I(\col_select_trans[4].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__C (.I(\col_select_trans[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06044__I (.I(\col_select_trans[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__A1 (.I(\col_select_trans[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A1 (.I(\col_select_trans[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06862__A1 (.I(\col_select_trans[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06043__I (.I(\col_select_trans[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(data_in_a[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(data_in_a[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(data_in_a[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(data_in_a[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(data_in_a[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(data_in_a[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(data_in_a[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(data_in_a[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(data_in_a[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(data_in_a[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(data_in_a[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(data_in_a[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(data_in_a[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(data_in_a[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(data_in_a[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(data_in_a[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12050__D (.I(\data_in_trans[0].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12070__D (.I(\data_in_trans[10].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__I (.I(\data_in_trans[10].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__I (.I(\data_in_trans[10].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__I (.I(\data_in_trans[10].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__I (.I(\data_in_trans[10].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12072__D (.I(\data_in_trans[11].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__I (.I(\data_in_trans[11].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__I (.I(\data_in_trans[11].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__I (.I(\data_in_trans[11].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__I (.I(\data_in_trans[11].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12074__D (.I(\data_in_trans[12].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__I (.I(\data_in_trans[12].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__I (.I(\data_in_trans[12].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__I (.I(\data_in_trans[12].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__I (.I(\data_in_trans[12].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12076__D (.I(\data_in_trans[13].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__I (.I(\data_in_trans[13].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__I (.I(\data_in_trans[13].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__I (.I(\data_in_trans[13].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__I (.I(\data_in_trans[13].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12078__D (.I(\data_in_trans[14].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__I (.I(\data_in_trans[14].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__I (.I(\data_in_trans[14].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__I (.I(\data_in_trans[14].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__I (.I(\data_in_trans[14].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12080__D (.I(\data_in_trans[15].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09761__I (.I(\data_in_trans[15].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__I (.I(\data_in_trans[15].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__I (.I(\data_in_trans[15].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__I (.I(\data_in_trans[15].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12052__D (.I(\data_in_trans[1].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__I (.I(\data_in_trans[1].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__I (.I(\data_in_trans[1].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12054__D (.I(\data_in_trans[2].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__I (.I(\data_in_trans[2].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08040__I (.I(\data_in_trans[2].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12056__D (.I(\data_in_trans[3].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__I (.I(\data_in_trans[3].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08044__I (.I(\data_in_trans[3].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12058__D (.I(\data_in_trans[4].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__I (.I(\data_in_trans[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08049__I (.I(\data_in_trans[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12060__D (.I(\data_in_trans[5].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__I (.I(\data_in_trans[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__I (.I(\data_in_trans[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12062__D (.I(\data_in_trans[6].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__I (.I(\data_in_trans[6].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__I (.I(\data_in_trans[6].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__I (.I(\data_in_trans[6].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__I (.I(\data_in_trans[6].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__I (.I(\data_in_trans[7].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__I (.I(\data_in_trans[7].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08314__I (.I(\data_in_trans[7].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__I (.I(\data_in_trans[7].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12066__D (.I(\data_in_trans[8].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__I (.I(\data_in_trans[8].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09037__I (.I(\data_in_trans[8].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__I (.I(\data_in_trans[8].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__I (.I(\data_in_trans[8].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12068__D (.I(\data_in_trans[9].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__I (.I(\data_in_trans[9].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__I (.I(\data_in_trans[9].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08325__I (.I(\data_in_trans[9].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__I (.I(\data_in_trans[9].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(inverter_select_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12092__D (.I(\inverter_select_trans.A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06034__A1 (.I(\inverter_select_trans.data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(mem_address_a[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(mem_address_a[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(mem_address_a[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(mem_address_a[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(mem_address_a[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(mem_address_a[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(mem_address_a[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(mem_address_a[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(mem_address_a[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(mem_address_a[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12006__D (.I(\mem_address_trans[0].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__A2 (.I(\mem_address_trans[0].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08099__I (.I(\mem_address_trans[0].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08021__I (.I(\mem_address_trans[0].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12008__D (.I(\mem_address_trans[1].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__A1 (.I(\mem_address_trans[1].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__I (.I(\mem_address_trans[1].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__I (.I(\mem_address_trans[1].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12010__D (.I(\mem_address_trans[2].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12012__D (.I(\mem_address_trans[3].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12014__D (.I(\mem_address_trans[4].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__I (.I(\mem_address_trans[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__I (.I(\mem_address_trans[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12016__D (.I(\mem_address_trans[5].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12018__D (.I(\mem_address_trans[6].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11873__A1 (.I(\mem_address_trans[6].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10837__I (.I(\mem_address_trans[6].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__I (.I(\mem_address_trans[6].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11873__A2 (.I(\mem_address_trans[7].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__I (.I(\mem_address_trans[7].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A4 (.I(\mem_address_trans[7].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12022__D (.I(\mem_address_trans[8].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12024__D (.I(\mem_address_trans[9].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(mem_write_n_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12086__D (.I(\mem_write_n_trans.A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(output_active_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold1_I (.I(\output_active_trans.data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(row_col_select_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12088__D (.I(\row_col_select_trans.A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05998__A2 (.I(\row_col_select_trans.data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05997__A2 (.I(\row_col_select_trans.data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__I (.I(\row_col_select_trans.data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(row_select_a[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(row_select_a[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(row_select_a[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(row_select_a[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(row_select_a[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(row_select_a[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12026__D (.I(\row_select_trans[0].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__A1 (.I(\row_select_trans[0].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__I (.I(\row_select_trans[0].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12028__D (.I(\row_select_trans[1].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12030__D (.I(\row_select_trans[2].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12032__D (.I(\row_select_trans[3].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__I (.I(\row_select_trans[3].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06504__I (.I(\row_select_trans[3].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__A2 (.I(\row_select_trans[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06521__A2 (.I(\row_select_trans[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__I (.I(\row_select_trans[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06507__A2 (.I(\row_select_trans[4].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12036__D (.I(\row_select_trans[5].A ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__A2 (.I(\row_select_trans[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__I (.I(\row_select_trans[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06513__A1 (.I(\row_select_trans[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06507__A1 (.I(\row_select_trans[5].data_sync ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A1 (.I(\u2.active_mem[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__B2 (.I(\u2.active_mem[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A1 (.I(\u2.active_mem[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__B2 (.I(\u2.active_mem[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__B2 (.I(\u2.active_mem[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__A1 (.I(\u2.active_mem[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A1 (.I(\u2.active_mem[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__B2 (.I(\u2.active_mem[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__A1 (.I(\u2.driver_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06021__A1 (.I(\u2.driver_mem[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__A1 (.I(\u2.driver_mem[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06015__A1 (.I(\u2.driver_mem[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06014__A1 (.I(\u2.driver_mem[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__A1 (.I(\u2.driver_mem[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__A1 (.I(\u2.driver_mem[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__I1 (.I(\u2.mem[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07831__B2 (.I(\u2.mem[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__I1 (.I(\u2.mem[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__B2 (.I(\u2.mem[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__I1 (.I(\u2.mem[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__B2 (.I(\u2.mem[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__I1 (.I(\u2.mem[10][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__B2 (.I(\u2.mem[10][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__I1 (.I(\u2.mem[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07357__B2 (.I(\u2.mem[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__I1 (.I(\u2.mem[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__B2 (.I(\u2.mem[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__I1 (.I(\u2.mem[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__B2 (.I(\u2.mem[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__I1 (.I(\u2.mem[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__B2 (.I(\u2.mem[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08603__I1 (.I(\u2.mem[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__B2 (.I(\u2.mem[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__I1 (.I(\u2.mem[11][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07979__B2 (.I(\u2.mem[11][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__I1 (.I(\u2.mem[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__B2 (.I(\u2.mem[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__I1 (.I(\u2.mem[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07482__B2 (.I(\u2.mem[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__I1 (.I(\u2.mem[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07708__B2 (.I(\u2.mem[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08637__I1 (.I(\u2.mem[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__B2 (.I(\u2.mem[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__I1 (.I(\u2.mem[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__B2 (.I(\u2.mem[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08642__I1 (.I(\u2.mem[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__B2 (.I(\u2.mem[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__I1 (.I(\u2.mem[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__B2 (.I(\u2.mem[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__I1 (.I(\u2.mem[12][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__B2 (.I(\u2.mem[12][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__I1 (.I(\u2.mem[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__B2 (.I(\u2.mem[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__I1 (.I(\u2.mem[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__B2 (.I(\u2.mem[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__I1 (.I(\u2.mem[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07339__B2 (.I(\u2.mem[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__I1 (.I(\u2.mem[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07418__B2 (.I(\u2.mem[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__I1 (.I(\u2.mem[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__B2 (.I(\u2.mem[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__I1 (.I(\u2.mem[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__B2 (.I(\u2.mem[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__I1 (.I(\u2.mem[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__B2 (.I(\u2.mem[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__I1 (.I(\u2.mem[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07655__B2 (.I(\u2.mem[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__I1 (.I(\u2.mem[144][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06633__A1 (.I(\u2.mem[144][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06167__A1 (.I(\u2.mem[144][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__I1 (.I(\u2.mem[144][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__A1 (.I(\u2.mem[144][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__A1 (.I(\u2.mem[144][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11110__I1 (.I(\u2.mem[144][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06741__A1 (.I(\u2.mem[144][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06294__A1 (.I(\u2.mem[144][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__I1 (.I(\u2.mem[144][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__C1 (.I(\u2.mem[144][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__A1 (.I(\u2.mem[144][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__I1 (.I(\u2.mem[144][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06820__A1 (.I(\u2.mem[144][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06365__A1 (.I(\u2.mem[144][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__I1 (.I(\u2.mem[144][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__A1 (.I(\u2.mem[144][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06400__A1 (.I(\u2.mem[144][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__I1 (.I(\u2.mem[145][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06598__C1 (.I(\u2.mem[145][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06140__A1 (.I(\u2.mem[145][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11122__I1 (.I(\u2.mem[145][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06689__A1 (.I(\u2.mem[145][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06229__A1 (.I(\u2.mem[145][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11124__I1 (.I(\u2.mem[145][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__C1 (.I(\u2.mem[145][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A1 (.I(\u2.mem[145][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__I1 (.I(\u2.mem[145][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06777__A1 (.I(\u2.mem[145][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__A1 (.I(\u2.mem[145][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11128__I1 (.I(\u2.mem[145][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__C1 (.I(\u2.mem[145][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__A1 (.I(\u2.mem[145][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__I1 (.I(\u2.mem[145][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__A1 (.I(\u2.mem[145][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__A1 (.I(\u2.mem[145][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11135__I1 (.I(\u2.mem[146][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__A1 (.I(\u2.mem[146][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06188__A1 (.I(\u2.mem[146][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__I1 (.I(\u2.mem[146][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__A1 (.I(\u2.mem[146][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__A1 (.I(\u2.mem[146][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__I1 (.I(\u2.mem[146][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06787__A1 (.I(\u2.mem[146][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06334__A1 (.I(\u2.mem[146][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__I1 (.I(\u2.mem[146][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__A1 (.I(\u2.mem[146][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06369__A1 (.I(\u2.mem[146][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__I1 (.I(\u2.mem[146][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06853__A1 (.I(\u2.mem[146][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__A1 (.I(\u2.mem[146][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11154__I1 (.I(\u2.mem[147][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__B2 (.I(\u2.mem[147][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__A1 (.I(\u2.mem[147][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11156__I1 (.I(\u2.mem[147][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__B2 (.I(\u2.mem[147][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06238__A1 (.I(\u2.mem[147][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__I1 (.I(\u2.mem[147][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__B2 (.I(\u2.mem[147][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__A1 (.I(\u2.mem[147][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11160__I1 (.I(\u2.mem[147][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__B2 (.I(\u2.mem[147][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06336__A1 (.I(\u2.mem[147][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__I1 (.I(\u2.mem[147][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__B2 (.I(\u2.mem[147][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__A1 (.I(\u2.mem[147][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__I1 (.I(\u2.mem[147][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__B2 (.I(\u2.mem[147][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06406__A1 (.I(\u2.mem[147][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__I1 (.I(\u2.mem[148][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__A1 (.I(\u2.mem[148][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__B2 (.I(\u2.mem[148][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__I1 (.I(\u2.mem[148][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__B2 (.I(\u2.mem[148][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__A1 (.I(\u2.mem[148][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__I1 (.I(\u2.mem[148][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__A1 (.I(\u2.mem[148][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06291__B2 (.I(\u2.mem[148][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__I1 (.I(\u2.mem[148][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06817__A1 (.I(\u2.mem[148][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__B2 (.I(\u2.mem[148][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11183__I1 (.I(\u2.mem[149][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__B2 (.I(\u2.mem[149][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06091__B2 (.I(\u2.mem[149][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__I1 (.I(\u2.mem[149][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06694__A1 (.I(\u2.mem[149][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06246__B2 (.I(\u2.mem[149][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__I1 (.I(\u2.mem[149][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__B2 (.I(\u2.mem[149][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__B2 (.I(\u2.mem[149][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11189__I1 (.I(\u2.mem[149][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__B2 (.I(\u2.mem[149][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06321__B2 (.I(\u2.mem[149][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__I1 (.I(\u2.mem[149][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__A1 (.I(\u2.mem[149][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__B2 (.I(\u2.mem[149][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11193__I1 (.I(\u2.mem[149][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__B2 (.I(\u2.mem[149][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__B2 (.I(\u2.mem[149][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__I1 (.I(\u2.mem[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07708__A1 (.I(\u2.mem[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08731__I1 (.I(\u2.mem[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__A1 (.I(\u2.mem[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__I1 (.I(\u2.mem[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__A1 (.I(\u2.mem[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__I1 (.I(\u2.mem[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__A1 (.I(\u2.mem[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08738__I1 (.I(\u2.mem[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__A1 (.I(\u2.mem[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__I1 (.I(\u2.mem[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__A1 (.I(\u2.mem[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__I1 (.I(\u2.mem[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__A1 (.I(\u2.mem[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__I1 (.I(\u2.mem[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__A1 (.I(\u2.mem[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__I1 (.I(\u2.mem[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__A1 (.I(\u2.mem[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__I1 (.I(\u2.mem[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__A1 (.I(\u2.mem[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__I1 (.I(\u2.mem[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07655__A1 (.I(\u2.mem[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__I1 (.I(\u2.mem[150][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__B2 (.I(\u2.mem[150][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__B2 (.I(\u2.mem[150][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__I1 (.I(\u2.mem[150][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__B2 (.I(\u2.mem[150][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__B2 (.I(\u2.mem[150][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11207__I1 (.I(\u2.mem[150][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__A1 (.I(\u2.mem[150][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__B2 (.I(\u2.mem[150][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__I1 (.I(\u2.mem[150][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A1 (.I(\u2.mem[150][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__B2 (.I(\u2.mem[150][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__I1 (.I(\u2.mem[150][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__B2 (.I(\u2.mem[150][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06344__B2 (.I(\u2.mem[150][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__I1 (.I(\u2.mem[150][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__A1 (.I(\u2.mem[150][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06379__B2 (.I(\u2.mem[150][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11223__I1 (.I(\u2.mem[151][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__A1 (.I(\u2.mem[151][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06071__B2 (.I(\u2.mem[151][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__I1 (.I(\u2.mem[151][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__A1 (.I(\u2.mem[151][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06231__B2 (.I(\u2.mem[151][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11227__I1 (.I(\u2.mem[151][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06738__A1 (.I(\u2.mem[151][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__B2 (.I(\u2.mem[151][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11229__I1 (.I(\u2.mem[151][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__A1 (.I(\u2.mem[151][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06317__B2 (.I(\u2.mem[151][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11231__I1 (.I(\u2.mem[151][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__A1 (.I(\u2.mem[151][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__B2 (.I(\u2.mem[151][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__I1 (.I(\u2.mem[151][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06841__A1 (.I(\u2.mem[151][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__B2 (.I(\u2.mem[151][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11238__I1 (.I(\u2.mem[152][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__B2 (.I(\u2.mem[152][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__A1 (.I(\u2.mem[152][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__I1 (.I(\u2.mem[152][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__B2 (.I(\u2.mem[152][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06291__A1 (.I(\u2.mem[152][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11244__I1 (.I(\u2.mem[152][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06767__B2 (.I(\u2.mem[152][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__A1 (.I(\u2.mem[152][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11248__I1 (.I(\u2.mem[152][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__B2 (.I(\u2.mem[152][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__A1 (.I(\u2.mem[152][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__I1 (.I(\u2.mem[153][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__A1 (.I(\u2.mem[153][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06204__A1 (.I(\u2.mem[153][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__I1 (.I(\u2.mem[153][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__A1 (.I(\u2.mem[153][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__B2 (.I(\u2.mem[153][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__I1 (.I(\u2.mem[153][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06745__A1 (.I(\u2.mem[153][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__A1 (.I(\u2.mem[153][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__I1 (.I(\u2.mem[153][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06765__A1 (.I(\u2.mem[153][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06327__A1 (.I(\u2.mem[153][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__I1 (.I(\u2.mem[153][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06846__A1 (.I(\u2.mem[153][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06396__A1 (.I(\u2.mem[153][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11267__I1 (.I(\u2.mem[154][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__A1 (.I(\u2.mem[154][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__A1 (.I(\u2.mem[154][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__I1 (.I(\u2.mem[154][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__A1 (.I(\u2.mem[154][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__B2 (.I(\u2.mem[154][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__I1 (.I(\u2.mem[154][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__A1 (.I(\u2.mem[154][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__A1 (.I(\u2.mem[154][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__I1 (.I(\u2.mem[154][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06763__A1 (.I(\u2.mem[154][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06330__A1 (.I(\u2.mem[154][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__I1 (.I(\u2.mem[154][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__A1 (.I(\u2.mem[154][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__A1 (.I(\u2.mem[154][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__I1 (.I(\u2.mem[155][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__A1 (.I(\u2.mem[155][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06155__B2 (.I(\u2.mem[155][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__I1 (.I(\u2.mem[155][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__A1 (.I(\u2.mem[155][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__B2 (.I(\u2.mem[155][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__I1 (.I(\u2.mem[155][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06728__A1 (.I(\u2.mem[155][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06277__B2 (.I(\u2.mem[155][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11292__I1 (.I(\u2.mem[155][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06780__A1 (.I(\u2.mem[155][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__A1 (.I(\u2.mem[155][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11294__I1 (.I(\u2.mem[155][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__A1 (.I(\u2.mem[155][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__B2 (.I(\u2.mem[155][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__I1 (.I(\u2.mem[155][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__A1 (.I(\u2.mem[155][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06378__B2 (.I(\u2.mem[155][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__I1 (.I(\u2.mem[156][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06664__B2 (.I(\u2.mem[156][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__B2 (.I(\u2.mem[156][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__I1 (.I(\u2.mem[156][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__B2 (.I(\u2.mem[156][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__B2 (.I(\u2.mem[156][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__I1 (.I(\u2.mem[156][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__B2 (.I(\u2.mem[156][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06296__B2 (.I(\u2.mem[156][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__I1 (.I(\u2.mem[156][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__B2 (.I(\u2.mem[156][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__B2 (.I(\u2.mem[156][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__I1 (.I(\u2.mem[156][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__B2 (.I(\u2.mem[156][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06367__B2 (.I(\u2.mem[156][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11315__I1 (.I(\u2.mem[157][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__B2 (.I(\u2.mem[157][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__B2 (.I(\u2.mem[157][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__I1 (.I(\u2.mem[157][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__B2 (.I(\u2.mem[157][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__B2 (.I(\u2.mem[157][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__I1 (.I(\u2.mem[157][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__B2 (.I(\u2.mem[157][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06266__B2 (.I(\u2.mem[157][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__I1 (.I(\u2.mem[157][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__B2 (.I(\u2.mem[157][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06308__B2 (.I(\u2.mem[157][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11323__I1 (.I(\u2.mem[157][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__B2 (.I(\u2.mem[157][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06348__B2 (.I(\u2.mem[157][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11330__I1 (.I(\u2.mem[158][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__B2 (.I(\u2.mem[158][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06071__A1 (.I(\u2.mem[158][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__I1 (.I(\u2.mem[158][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__B2 (.I(\u2.mem[158][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06231__A1 (.I(\u2.mem[158][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__I1 (.I(\u2.mem[158][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06738__B2 (.I(\u2.mem[158][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__A1 (.I(\u2.mem[158][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__I1 (.I(\u2.mem[158][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__B2 (.I(\u2.mem[158][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06317__A1 (.I(\u2.mem[158][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11342__I1 (.I(\u2.mem[158][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__B2 (.I(\u2.mem[158][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__A1 (.I(\u2.mem[158][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__I1 (.I(\u2.mem[158][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06841__B2 (.I(\u2.mem[158][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__A1 (.I(\u2.mem[158][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__I1 (.I(\u2.mem[159][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__A1 (.I(\u2.mem[159][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06098__B2 (.I(\u2.mem[159][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11351__I1 (.I(\u2.mem[159][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__C1 (.I(\u2.mem[159][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06246__A1 (.I(\u2.mem[159][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__I1 (.I(\u2.mem[159][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__A1 (.I(\u2.mem[159][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__A1 (.I(\u2.mem[159][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__I1 (.I(\u2.mem[159][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__A1 (.I(\u2.mem[159][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06321__A1 (.I(\u2.mem[159][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11357__I1 (.I(\u2.mem[159][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__C1 (.I(\u2.mem[159][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__A1 (.I(\u2.mem[159][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__I1 (.I(\u2.mem[159][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__A1 (.I(\u2.mem[159][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__A1 (.I(\u2.mem[159][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11365__I1 (.I(\u2.mem[160][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__B2 (.I(\u2.mem[160][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06204__B2 (.I(\u2.mem[160][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__I1 (.I(\u2.mem[160][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06745__B2 (.I(\u2.mem[160][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__B2 (.I(\u2.mem[160][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11371__I1 (.I(\u2.mem[160][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06765__B2 (.I(\u2.mem[160][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06327__B2 (.I(\u2.mem[160][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__I1 (.I(\u2.mem[161][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__B2 (.I(\u2.mem[161][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06091__C2 (.I(\u2.mem[161][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11381__I1 (.I(\u2.mem[161][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__B2 (.I(\u2.mem[161][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06249__B2 (.I(\u2.mem[161][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11383__I1 (.I(\u2.mem[161][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__B2 (.I(\u2.mem[161][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__B2 (.I(\u2.mem[161][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__I1 (.I(\u2.mem[161][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__B2 (.I(\u2.mem[161][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06323__B2 (.I(\u2.mem[161][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__I1 (.I(\u2.mem[161][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__B2 (.I(\u2.mem[161][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__B2 (.I(\u2.mem[161][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11389__I1 (.I(\u2.mem[161][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__B2 (.I(\u2.mem[161][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__B2 (.I(\u2.mem[161][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__I1 (.I(\u2.mem[162][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__B2 (.I(\u2.mem[162][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__B2 (.I(\u2.mem[162][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__I1 (.I(\u2.mem[162][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__C2 (.I(\u2.mem[162][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__C1 (.I(\u2.mem[162][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11400__I1 (.I(\u2.mem[162][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__B2 (.I(\u2.mem[162][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__B2 (.I(\u2.mem[162][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__I1 (.I(\u2.mem[162][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06763__B2 (.I(\u2.mem[162][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06330__B2 (.I(\u2.mem[162][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11406__I1 (.I(\u2.mem[162][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__B2 (.I(\u2.mem[162][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__B2 (.I(\u2.mem[162][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__I1 (.I(\u2.mem[162][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06849__B2 (.I(\u2.mem[162][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__B2 (.I(\u2.mem[162][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__I1 (.I(\u2.mem[163][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06598__B2 (.I(\u2.mem[163][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06140__B2 (.I(\u2.mem[163][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__I1 (.I(\u2.mem[163][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06705__B2 (.I(\u2.mem[163][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06224__A1 (.I(\u2.mem[163][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__I1 (.I(\u2.mem[163][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__B2 (.I(\u2.mem[163][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__B2 (.I(\u2.mem[163][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__I1 (.I(\u2.mem[163][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__B2 (.I(\u2.mem[163][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__C1 (.I(\u2.mem[163][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__I1 (.I(\u2.mem[163][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__B2 (.I(\u2.mem[163][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__B2 (.I(\u2.mem[163][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11423__I1 (.I(\u2.mem[163][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__B2 (.I(\u2.mem[163][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__C1 (.I(\u2.mem[163][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11428__I1 (.I(\u2.mem[164][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A1 (.I(\u2.mem[164][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06114__B2 (.I(\u2.mem[164][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11430__I1 (.I(\u2.mem[164][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06696__A1 (.I(\u2.mem[164][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__B2 (.I(\u2.mem[164][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11432__I1 (.I(\u2.mem[164][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__A1 (.I(\u2.mem[164][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__B2 (.I(\u2.mem[164][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__I1 (.I(\u2.mem[164][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__A1 (.I(\u2.mem[164][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06306__B2 (.I(\u2.mem[164][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11436__I1 (.I(\u2.mem[164][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06797__A1 (.I(\u2.mem[164][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06346__B2 (.I(\u2.mem[164][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11438__I1 (.I(\u2.mem[164][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06826__A1 (.I(\u2.mem[164][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06381__B2 (.I(\u2.mem[164][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__I1 (.I(\u2.mem[165][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06598__A1 (.I(\u2.mem[165][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06140__C1 (.I(\u2.mem[165][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11444__I1 (.I(\u2.mem[165][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06705__A1 (.I(\u2.mem[165][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06224__B2 (.I(\u2.mem[165][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11446__I1 (.I(\u2.mem[165][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__A1 (.I(\u2.mem[165][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__C1 (.I(\u2.mem[165][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__I1 (.I(\u2.mem[165][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__A1 (.I(\u2.mem[165][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__B2 (.I(\u2.mem[165][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11450__I1 (.I(\u2.mem[165][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__A1 (.I(\u2.mem[165][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__C1 (.I(\u2.mem[165][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__I1 (.I(\u2.mem[165][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__A1 (.I(\u2.mem[165][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__B2 (.I(\u2.mem[165][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11478__I1 (.I(\u2.mem[166][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__A1 (.I(\u2.mem[166][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__A1 (.I(\u2.mem[166][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__I1 (.I(\u2.mem[167][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06578__A1 (.I(\u2.mem[167][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__A1 (.I(\u2.mem[167][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11484__I1 (.I(\u2.mem[167][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06697__A1 (.I(\u2.mem[167][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06241__A1 (.I(\u2.mem[167][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11486__I1 (.I(\u2.mem[167][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__A1 (.I(\u2.mem[167][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__A1 (.I(\u2.mem[167][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__I1 (.I(\u2.mem[167][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06770__A1 (.I(\u2.mem[167][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__A1 (.I(\u2.mem[167][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11497__I1 (.I(\u2.mem[168][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06610__B2 (.I(\u2.mem[168][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06083__B2 (.I(\u2.mem[168][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11503__I1 (.I(\u2.mem[168][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06774__A1 (.I(\u2.mem[168][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__B2 (.I(\u2.mem[168][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11505__I1 (.I(\u2.mem[168][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__C1 (.I(\u2.mem[168][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__C2 (.I(\u2.mem[168][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11507__I1 (.I(\u2.mem[168][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__B2 (.I(\u2.mem[168][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__B2 (.I(\u2.mem[168][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11511__I1 (.I(\u2.mem[169][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__A1 (.I(\u2.mem[169][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__B2 (.I(\u2.mem[169][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__I1 (.I(\u2.mem[169][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__A1 (.I(\u2.mem[169][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__B2 (.I(\u2.mem[169][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11519__I1 (.I(\u2.mem[169][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__A1 (.I(\u2.mem[169][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__B2 (.I(\u2.mem[169][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__I1 (.I(\u2.mem[16][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__A1 (.I(\u2.mem[16][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11526__I1 (.I(\u2.mem[170][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06664__A1 (.I(\u2.mem[170][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__A1 (.I(\u2.mem[170][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11529__I1 (.I(\u2.mem[170][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__A1 (.I(\u2.mem[170][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__A1 (.I(\u2.mem[170][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11532__I1 (.I(\u2.mem[170][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__A1 (.I(\u2.mem[170][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06296__A1 (.I(\u2.mem[170][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__I1 (.I(\u2.mem[170][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__A1 (.I(\u2.mem[170][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__A1 (.I(\u2.mem[170][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11545__I1 (.I(\u2.mem[171][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__A1 (.I(\u2.mem[171][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__A1 (.I(\u2.mem[171][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11547__I1 (.I(\u2.mem[171][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__A1 (.I(\u2.mem[171][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__A1 (.I(\u2.mem[171][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11549__I1 (.I(\u2.mem[171][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__A1 (.I(\u2.mem[171][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06266__A1 (.I(\u2.mem[171][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__I1 (.I(\u2.mem[171][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__A1 (.I(\u2.mem[171][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06308__A1 (.I(\u2.mem[171][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11553__I1 (.I(\u2.mem[171][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__A1 (.I(\u2.mem[171][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06348__A1 (.I(\u2.mem[171][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11555__I1 (.I(\u2.mem[171][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__A1 (.I(\u2.mem[171][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__A1 (.I(\u2.mem[171][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11560__I1 (.I(\u2.mem[172][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06536__B2 (.I(\u2.mem[172][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__C1 (.I(\u2.mem[172][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11562__I1 (.I(\u2.mem[172][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__B2 (.I(\u2.mem[172][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__C1 (.I(\u2.mem[172][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11566__I1 (.I(\u2.mem[172][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06779__B2 (.I(\u2.mem[172][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__A1 (.I(\u2.mem[172][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11568__I1 (.I(\u2.mem[172][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__B2 (.I(\u2.mem[172][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06344__A1 (.I(\u2.mem[172][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11570__I1 (.I(\u2.mem[172][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06833__B2 (.I(\u2.mem[172][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06377__C1 (.I(\u2.mem[172][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11574__I1 (.I(\u2.mem[173][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06639__B2 (.I(\u2.mem[173][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__A1 (.I(\u2.mem[173][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11576__I1 (.I(\u2.mem[173][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06682__B2 (.I(\u2.mem[173][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06233__A1 (.I(\u2.mem[173][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__I1 (.I(\u2.mem[173][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06787__B2 (.I(\u2.mem[173][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06331__A1 (.I(\u2.mem[173][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11589__I1 (.I(\u2.mem[174][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__B2 (.I(\u2.mem[174][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06155__A1 (.I(\u2.mem[174][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11592__I1 (.I(\u2.mem[174][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__B2 (.I(\u2.mem[174][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__A1 (.I(\u2.mem[174][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11598__I1 (.I(\u2.mem[174][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__B2 (.I(\u2.mem[174][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__A1 (.I(\u2.mem[174][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11601__I1 (.I(\u2.mem[174][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__A1 (.I(\u2.mem[174][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__A1 (.I(\u2.mem[174][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11608__I1 (.I(\u2.mem[175][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__B2 (.I(\u2.mem[175][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06098__A1 (.I(\u2.mem[175][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11616__I1 (.I(\u2.mem[175][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__B2 (.I(\u2.mem[175][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__A1 (.I(\u2.mem[175][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11624__I1 (.I(\u2.mem[176][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06536__A1 (.I(\u2.mem[176][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__B2 (.I(\u2.mem[176][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__I1 (.I(\u2.mem[176][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__A1 (.I(\u2.mem[176][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__B2 (.I(\u2.mem[176][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11628__I1 (.I(\u2.mem[176][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06729__A1 (.I(\u2.mem[176][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__C2 (.I(\u2.mem[176][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11638__I1 (.I(\u2.mem[177][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06610__A1 (.I(\u2.mem[177][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06083__A1 (.I(\u2.mem[177][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__I1 (.I(\u2.mem[177][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06705__C2 (.I(\u2.mem[177][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06229__B2 (.I(\u2.mem[177][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__I1 (.I(\u2.mem[177][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06739__A1 (.I(\u2.mem[177][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06287__B2 (.I(\u2.mem[177][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11653__I1 (.I(\u2.mem[178][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__B2 (.I(\u2.mem[178][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06114__A1 (.I(\u2.mem[178][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11656__I1 (.I(\u2.mem[178][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06696__B2 (.I(\u2.mem[178][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__A1 (.I(\u2.mem[178][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11659__I1 (.I(\u2.mem[178][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__B2 (.I(\u2.mem[178][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A1 (.I(\u2.mem[178][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11662__I1 (.I(\u2.mem[178][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__B2 (.I(\u2.mem[178][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06306__A1 (.I(\u2.mem[178][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11665__I1 (.I(\u2.mem[178][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06797__B2 (.I(\u2.mem[178][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06346__A1 (.I(\u2.mem[178][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11672__I1 (.I(\u2.mem[179][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06669__A1 (.I(\u2.mem[179][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__B2 (.I(\u2.mem[179][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11674__I1 (.I(\u2.mem[179][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06684__A1 (.I(\u2.mem[179][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06235__B2 (.I(\u2.mem[179][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11676__I1 (.I(\u2.mem[179][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__A1 (.I(\u2.mem[179][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__B2 (.I(\u2.mem[179][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11678__I1 (.I(\u2.mem[179][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06785__A1 (.I(\u2.mem[179][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06333__B2 (.I(\u2.mem[179][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11680__I1 (.I(\u2.mem[179][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__A1 (.I(\u2.mem[179][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__B2 (.I(\u2.mem[179][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11687__I1 (.I(\u2.mem[180][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__A1 (.I(\u2.mem[180][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__A1 (.I(\u2.mem[180][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11689__I1 (.I(\u2.mem[180][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__A1 (.I(\u2.mem[180][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__A1 (.I(\u2.mem[180][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11691__I1 (.I(\u2.mem[180][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06730__A1 (.I(\u2.mem[180][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__B2 (.I(\u2.mem[180][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11693__I1 (.I(\u2.mem[180][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06779__A1 (.I(\u2.mem[180][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__B2 (.I(\u2.mem[180][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11695__I1 (.I(\u2.mem[180][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__A1 (.I(\u2.mem[180][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__B2 (.I(\u2.mem[180][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11697__I1 (.I(\u2.mem[180][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06833__A1 (.I(\u2.mem[180][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06379__A1 (.I(\u2.mem[180][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11701__I1 (.I(\u2.mem[181][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__C1 (.I(\u2.mem[181][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06155__C2 (.I(\u2.mem[181][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11703__I1 (.I(\u2.mem[181][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__C1 (.I(\u2.mem[181][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__C2 (.I(\u2.mem[181][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11705__I1 (.I(\u2.mem[181][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06728__C1 (.I(\u2.mem[181][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06277__C2 (.I(\u2.mem[181][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11707__I1 (.I(\u2.mem[181][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__C1 (.I(\u2.mem[181][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__C2 (.I(\u2.mem[181][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11709__I1 (.I(\u2.mem[181][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__B2 (.I(\u2.mem[181][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__C2 (.I(\u2.mem[181][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11711__I1 (.I(\u2.mem[181][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__C1 (.I(\u2.mem[181][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06378__C2 (.I(\u2.mem[181][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11716__I1 (.I(\u2.mem[182][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06633__B2 (.I(\u2.mem[182][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06167__B2 (.I(\u2.mem[182][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11719__I1 (.I(\u2.mem[182][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__B2 (.I(\u2.mem[182][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__B2 (.I(\u2.mem[182][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11722__I1 (.I(\u2.mem[182][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06741__B2 (.I(\u2.mem[182][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06294__B2 (.I(\u2.mem[182][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11725__I1 (.I(\u2.mem[182][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__B2 (.I(\u2.mem[182][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__B2 (.I(\u2.mem[182][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11731__I1 (.I(\u2.mem[182][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__B2 (.I(\u2.mem[182][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06400__B2 (.I(\u2.mem[182][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11735__I1 (.I(\u2.mem[183][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06578__B2 (.I(\u2.mem[183][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__B2 (.I(\u2.mem[183][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11737__I1 (.I(\u2.mem[183][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06697__B2 (.I(\u2.mem[183][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06241__B2 (.I(\u2.mem[183][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11739__I1 (.I(\u2.mem[183][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__B2 (.I(\u2.mem[183][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__B2 (.I(\u2.mem[183][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11741__I1 (.I(\u2.mem[183][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06770__B2 (.I(\u2.mem[183][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__B2 (.I(\u2.mem[183][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11743__I1 (.I(\u2.mem[183][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06798__B2 (.I(\u2.mem[183][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06347__B2 (.I(\u2.mem[183][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11745__I1 (.I(\u2.mem[183][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06827__B2 (.I(\u2.mem[183][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__B2 (.I(\u2.mem[183][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11750__I1 (.I(\u2.mem[184][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__A1 (.I(\u2.mem[184][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__A1 (.I(\u2.mem[184][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11752__I1 (.I(\u2.mem[184][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06698__A1 (.I(\u2.mem[184][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06244__A1 (.I(\u2.mem[184][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11754__I1 (.I(\u2.mem[184][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__A1 (.I(\u2.mem[184][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06274__A1 (.I(\u2.mem[184][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11756__I1 (.I(\u2.mem[184][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06772__A1 (.I(\u2.mem[184][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06309__A1 (.I(\u2.mem[184][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11758__I1 (.I(\u2.mem[184][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__A1 (.I(\u2.mem[184][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06349__A1 (.I(\u2.mem[184][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11760__I1 (.I(\u2.mem[184][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06828__A1 (.I(\u2.mem[184][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06384__A1 (.I(\u2.mem[184][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11764__I1 (.I(\u2.mem[185][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06639__A1 (.I(\u2.mem[185][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__B2 (.I(\u2.mem[185][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11766__I1 (.I(\u2.mem[185][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06682__A1 (.I(\u2.mem[185][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06233__B2 (.I(\u2.mem[185][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11768__I1 (.I(\u2.mem[185][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06749__A1 (.I(\u2.mem[185][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__B2 (.I(\u2.mem[185][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11770__I1 (.I(\u2.mem[185][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__A1 (.I(\u2.mem[185][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06331__B2 (.I(\u2.mem[185][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11772__I1 (.I(\u2.mem[185][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__A1 (.I(\u2.mem[185][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__B2 (.I(\u2.mem[185][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11774__I1 (.I(\u2.mem[185][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__A1 (.I(\u2.mem[185][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__B2 (.I(\u2.mem[185][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11779__I1 (.I(\u2.mem[186][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__B2 (.I(\u2.mem[186][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06188__B2 (.I(\u2.mem[186][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11788__I1 (.I(\u2.mem[186][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__C2 (.I(\u2.mem[186][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06334__B2 (.I(\u2.mem[186][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11791__I1 (.I(\u2.mem[186][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__B2 (.I(\u2.mem[186][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06369__B2 (.I(\u2.mem[186][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11794__I1 (.I(\u2.mem[186][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06853__B2 (.I(\u2.mem[186][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__B2 (.I(\u2.mem[186][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11798__I1 (.I(\u2.mem[187][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__A1 (.I(\u2.mem[187][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06130__B2 (.I(\u2.mem[187][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11800__I1 (.I(\u2.mem[187][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__B2 (.I(\u2.mem[187][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06250__A1 (.I(\u2.mem[187][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11802__I1 (.I(\u2.mem[187][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06732__A1 (.I(\u2.mem[187][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06280__A1 (.I(\u2.mem[187][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11804__I1 (.I(\u2.mem[187][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__A1 (.I(\u2.mem[187][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A1 (.I(\u2.mem[187][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11806__I1 (.I(\u2.mem[187][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06802__B2 (.I(\u2.mem[187][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__A1 (.I(\u2.mem[187][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11808__I1 (.I(\u2.mem[187][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06835__A1 (.I(\u2.mem[187][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06389__A1 (.I(\u2.mem[187][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11813__I1 (.I(\u2.mem[188][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__A1 (.I(\u2.mem[188][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06130__A1 (.I(\u2.mem[188][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11815__I1 (.I(\u2.mem[188][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__A1 (.I(\u2.mem[188][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__B2 (.I(\u2.mem[188][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11817__I1 (.I(\u2.mem[188][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06733__A1 (.I(\u2.mem[188][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__B2 (.I(\u2.mem[188][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11819__I1 (.I(\u2.mem[188][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06760__A1 (.I(\u2.mem[188][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__B2 (.I(\u2.mem[188][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11821__I1 (.I(\u2.mem[188][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06802__A1 (.I(\u2.mem[188][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__B2 (.I(\u2.mem[188][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11823__I1 (.I(\u2.mem[188][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__A1 (.I(\u2.mem[188][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__B2 (.I(\u2.mem[188][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11827__I1 (.I(\u2.mem[189][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06536__C2 (.I(\u2.mem[189][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__A1 (.I(\u2.mem[189][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11829__I1 (.I(\u2.mem[189][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__C2 (.I(\u2.mem[189][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__A1 (.I(\u2.mem[189][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11831__I1 (.I(\u2.mem[189][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06729__B2 (.I(\u2.mem[189][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__A1 (.I(\u2.mem[189][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11833__I1 (.I(\u2.mem[189][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__B2 (.I(\u2.mem[189][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06313__A1 (.I(\u2.mem[189][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11835__I1 (.I(\u2.mem[189][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__B2 (.I(\u2.mem[189][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__A1 (.I(\u2.mem[189][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11837__I1 (.I(\u2.mem[189][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06832__B2 (.I(\u2.mem[189][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06377__A1 (.I(\u2.mem[189][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__I1 (.I(\u2.mem[18][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A1 (.I(\u2.mem[18][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11842__I1 (.I(\u2.mem[190][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__B2 (.I(\u2.mem[190][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06199__A1 (.I(\u2.mem[190][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11845__I1 (.I(\u2.mem[190][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06717__B2 (.I(\u2.mem[190][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06257__A1 (.I(\u2.mem[190][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11848__I1 (.I(\u2.mem[190][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06744__B2 (.I(\u2.mem[190][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06289__A1 (.I(\u2.mem[190][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11851__I1 (.I(\u2.mem[190][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__B2 (.I(\u2.mem[190][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06326__A1 (.I(\u2.mem[190][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11854__I1 (.I(\u2.mem[190][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__B2 (.I(\u2.mem[190][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06360__A1 (.I(\u2.mem[190][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11857__I1 (.I(\u2.mem[190][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__B2 (.I(\u2.mem[190][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__A1 (.I(\u2.mem[190][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11861__I1 (.I(\u2.mem[191][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06669__B2 (.I(\u2.mem[191][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__A1 (.I(\u2.mem[191][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11863__I1 (.I(\u2.mem[191][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06684__B2 (.I(\u2.mem[191][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06235__A1 (.I(\u2.mem[191][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11865__I1 (.I(\u2.mem[191][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__B2 (.I(\u2.mem[191][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__A1 (.I(\u2.mem[191][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11867__I1 (.I(\u2.mem[191][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06785__B2 (.I(\u2.mem[191][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06333__A1 (.I(\u2.mem[191][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11869__I1 (.I(\u2.mem[191][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__B2 (.I(\u2.mem[191][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__A1 (.I(\u2.mem[191][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11871__I1 (.I(\u2.mem[191][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06852__B2 (.I(\u2.mem[191][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__A1 (.I(\u2.mem[191][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11878__I0 (.I(\u2.mem[192][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__B2 (.I(\u2.mem[192][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__B2 (.I(\u2.mem[192][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06130__C2 (.I(\u2.mem[192][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11880__I0 (.I(\u2.mem[192][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__C2 (.I(\u2.mem[192][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__B2 (.I(\u2.mem[192][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06250__B2 (.I(\u2.mem[192][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11883__I0 (.I(\u2.mem[192][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06732__B2 (.I(\u2.mem[192][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06433__A1 (.I(\u2.mem[192][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06280__B2 (.I(\u2.mem[192][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11885__I0 (.I(\u2.mem[192][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__B2 (.I(\u2.mem[192][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__A1 (.I(\u2.mem[192][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__B2 (.I(\u2.mem[192][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11887__I0 (.I(\u2.mem[192][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06802__C2 (.I(\u2.mem[192][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__B2 (.I(\u2.mem[192][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__B2 (.I(\u2.mem[192][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11889__I0 (.I(\u2.mem[192][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06835__B2 (.I(\u2.mem[192][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06445__A1 (.I(\u2.mem[192][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06389__B2 (.I(\u2.mem[192][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11915__I1 (.I(\u2.mem[193][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__C1 (.I(\u2.mem[193][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__A1 (.I(\u2.mem[193][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06071__C2 (.I(\u2.mem[193][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11937__I1 (.I(\u2.mem[193][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__A1 (.I(\u2.mem[193][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11939__I1 (.I(\u2.mem[193][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__A1 (.I(\u2.mem[193][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11917__I1 (.I(\u2.mem[193][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__C1 (.I(\u2.mem[193][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__A1 (.I(\u2.mem[193][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A1 (.I(\u2.mem[193][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11919__I1 (.I(\u2.mem[193][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06739__B2 (.I(\u2.mem[193][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06436__A1 (.I(\u2.mem[193][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06287__A1 (.I(\u2.mem[193][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11921__I1 (.I(\u2.mem[193][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__C1 (.I(\u2.mem[193][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__A1 (.I(\u2.mem[193][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06317__C2 (.I(\u2.mem[193][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11924__I1 (.I(\u2.mem[193][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__B2 (.I(\u2.mem[193][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__A1 (.I(\u2.mem[193][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06353__A1 (.I(\u2.mem[193][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11926__I1 (.I(\u2.mem[193][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06841__C1 (.I(\u2.mem[193][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__A1 (.I(\u2.mem[193][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__C2 (.I(\u2.mem[193][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11933__I1 (.I(\u2.mem[193][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__A1 (.I(\u2.mem[193][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11935__I1 (.I(\u2.mem[193][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__A1 (.I(\u2.mem[193][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11953__I1 (.I(\u2.mem[194][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__A1 (.I(\u2.mem[194][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__A1 (.I(\u2.mem[194][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06199__B2 (.I(\u2.mem[194][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11955__I1 (.I(\u2.mem[194][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06717__A1 (.I(\u2.mem[194][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__A1 (.I(\u2.mem[194][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06257__C2 (.I(\u2.mem[194][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11958__I1 (.I(\u2.mem[194][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06744__A1 (.I(\u2.mem[194][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06436__B2 (.I(\u2.mem[194][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06289__B2 (.I(\u2.mem[194][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11960__I1 (.I(\u2.mem[194][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__A1 (.I(\u2.mem[194][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__B2 (.I(\u2.mem[194][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06326__B2 (.I(\u2.mem[194][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11962__I1 (.I(\u2.mem[194][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__A1 (.I(\u2.mem[194][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__A1 (.I(\u2.mem[194][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06360__B2 (.I(\u2.mem[194][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11964__I1 (.I(\u2.mem[194][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__A1 (.I(\u2.mem[194][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__B2 (.I(\u2.mem[194][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__B2 (.I(\u2.mem[194][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11971__I1 (.I(\u2.mem[194][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__B2 (.I(\u2.mem[194][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11973__I1 (.I(\u2.mem[194][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__B2 (.I(\u2.mem[194][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__I1 (.I(\u2.mem[19][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__B2 (.I(\u2.mem[19][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__I1 (.I(\u2.mem[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07377__B2 (.I(\u2.mem[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__I1 (.I(\u2.mem[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__B2 (.I(\u2.mem[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__I1 (.I(\u2.mem[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__B2 (.I(\u2.mem[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__I1 (.I(\u2.mem[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__A1 (.I(\u2.mem[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__I1 (.I(\u2.mem[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__B2 (.I(\u2.mem[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__I1 (.I(\u2.mem[20][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__B2 (.I(\u2.mem[20][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__I1 (.I(\u2.mem[20][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__B2 (.I(\u2.mem[20][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__I1 (.I(\u2.mem[20][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07817__B2 (.I(\u2.mem[20][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__I1 (.I(\u2.mem[20][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__B2 (.I(\u2.mem[20][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__I1 (.I(\u2.mem[20][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__B2 (.I(\u2.mem[20][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__I1 (.I(\u2.mem[20][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07970__B2 (.I(\u2.mem[20][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__I1 (.I(\u2.mem[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__B2 (.I(\u2.mem[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__I1 (.I(\u2.mem[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__B2 (.I(\u2.mem[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__I1 (.I(\u2.mem[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__B2 (.I(\u2.mem[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__I1 (.I(\u2.mem[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07343__B2 (.I(\u2.mem[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__I1 (.I(\u2.mem[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07422__B2 (.I(\u2.mem[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__I1 (.I(\u2.mem[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__B2 (.I(\u2.mem[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__I1 (.I(\u2.mem[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__B2 (.I(\u2.mem[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__I1 (.I(\u2.mem[20][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__B2 (.I(\u2.mem[20][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__I1 (.I(\u2.mem[20][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__B2 (.I(\u2.mem[20][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__I1 (.I(\u2.mem[21][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__B2 (.I(\u2.mem[21][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__I1 (.I(\u2.mem[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07374__B2 (.I(\u2.mem[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__I1 (.I(\u2.mem[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07443__B2 (.I(\u2.mem[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__I1 (.I(\u2.mem[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__B2 (.I(\u2.mem[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__I1 (.I(\u2.mem[22][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__B2 (.I(\u2.mem[22][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__I1 (.I(\u2.mem[22][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__B2 (.I(\u2.mem[22][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__I1 (.I(\u2.mem[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__B2 (.I(\u2.mem[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__I1 (.I(\u2.mem[23][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__A1 (.I(\u2.mem[23][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__I1 (.I(\u2.mem[24][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__B2 (.I(\u2.mem[24][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__I1 (.I(\u2.mem[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07487__B2 (.I(\u2.mem[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__I1 (.I(\u2.mem[24][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__B2 (.I(\u2.mem[24][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__I1 (.I(\u2.mem[25][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07720__B2 (.I(\u2.mem[25][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__I1 (.I(\u2.mem[25][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__B2 (.I(\u2.mem[25][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09241__I1 (.I(\u2.mem[25][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__B2 (.I(\u2.mem[25][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__I1 (.I(\u2.mem[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__B2 (.I(\u2.mem[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09206__I1 (.I(\u2.mem[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07363__B2 (.I(\u2.mem[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09209__I1 (.I(\u2.mem[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__B2 (.I(\u2.mem[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__I1 (.I(\u2.mem[25][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07673__B2 (.I(\u2.mem[25][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09269__I1 (.I(\u2.mem[26][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07718__A1 (.I(\u2.mem[26][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__I1 (.I(\u2.mem[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07197__A1 (.I(\u2.mem[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09251__I1 (.I(\u2.mem[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07244__A1 (.I(\u2.mem[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__I1 (.I(\u2.mem[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__A1 (.I(\u2.mem[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09267__I1 (.I(\u2.mem[26][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__A1 (.I(\u2.mem[26][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__I1 (.I(\u2.mem[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__A1 (.I(\u2.mem[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__I1 (.I(\u2.mem[27][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A1 (.I(\u2.mem[27][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09313__I1 (.I(\u2.mem[27][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__A1 (.I(\u2.mem[27][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__I1 (.I(\u2.mem[27][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07869__A1 (.I(\u2.mem[27][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__I1 (.I(\u2.mem[27][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__A1 (.I(\u2.mem[27][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__I1 (.I(\u2.mem[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07160__A1 (.I(\u2.mem[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09290__I1 (.I(\u2.mem[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__A1 (.I(\u2.mem[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__I1 (.I(\u2.mem[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__A1 (.I(\u2.mem[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__I1 (.I(\u2.mem[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07315__A1 (.I(\u2.mem[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__I1 (.I(\u2.mem[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07397__A1 (.I(\u2.mem[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__I1 (.I(\u2.mem[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__A1 (.I(\u2.mem[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09301__I1 (.I(\u2.mem[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__A1 (.I(\u2.mem[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__I1 (.I(\u2.mem[27][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07552__A1 (.I(\u2.mem[27][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__I1 (.I(\u2.mem[27][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A1 (.I(\u2.mem[27][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__I1 (.I(\u2.mem[28][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__A1 (.I(\u2.mem[28][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__I1 (.I(\u2.mem[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__A1 (.I(\u2.mem[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__I1 (.I(\u2.mem[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__A1 (.I(\u2.mem[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09334__I1 (.I(\u2.mem[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07366__A1 (.I(\u2.mem[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__I1 (.I(\u2.mem[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__A1 (.I(\u2.mem[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__I1 (.I(\u2.mem[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07092__A1 (.I(\u2.mem[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__I1 (.I(\u2.mem[29][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__A1 (.I(\u2.mem[29][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__I1 (.I(\u2.mem[29][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__A1 (.I(\u2.mem[29][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__I1 (.I(\u2.mem[29][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__A1 (.I(\u2.mem[29][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__I1 (.I(\u2.mem[29][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07979__A1 (.I(\u2.mem[29][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__I1 (.I(\u2.mem[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__A1 (.I(\u2.mem[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__I1 (.I(\u2.mem[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__A1 (.I(\u2.mem[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09372__I1 (.I(\u2.mem[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07289__A1 (.I(\u2.mem[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09392__I1 (.I(\u2.mem[29][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__A1 (.I(\u2.mem[29][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__I1 (.I(\u2.mem[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06918__B2 (.I(\u2.mem[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08182__I1 (.I(\u2.mem[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__B2 (.I(\u2.mem[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__I1 (.I(\u2.mem[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07158__B2 (.I(\u2.mem[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__I1 (.I(\u2.mem[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__B2 (.I(\u2.mem[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__I1 (.I(\u2.mem[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__B2 (.I(\u2.mem[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__I1 (.I(\u2.mem[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__B2 (.I(\u2.mem[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09439__I1 (.I(\u2.mem[30][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__B2 (.I(\u2.mem[30][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__I1 (.I(\u2.mem[30][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__B2 (.I(\u2.mem[30][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__I1 (.I(\u2.mem[30][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__B2 (.I(\u2.mem[30][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09446__I1 (.I(\u2.mem[30][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__B2 (.I(\u2.mem[30][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__I1 (.I(\u2.mem[30][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__B2 (.I(\u2.mem[30][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__I1 (.I(\u2.mem[30][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07954__B2 (.I(\u2.mem[30][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__I1 (.I(\u2.mem[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07159__B2 (.I(\u2.mem[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__I1 (.I(\u2.mem[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07220__B2 (.I(\u2.mem[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__I1 (.I(\u2.mem[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__B2 (.I(\u2.mem[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__I1 (.I(\u2.mem[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__B2 (.I(\u2.mem[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__I1 (.I(\u2.mem[30][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__B2 (.I(\u2.mem[30][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__I1 (.I(\u2.mem[30][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07633__B2 (.I(\u2.mem[30][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__I1 (.I(\u2.mem[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__B2 (.I(\u2.mem[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__I1 (.I(\u2.mem[31][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__B2 (.I(\u2.mem[31][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__I1 (.I(\u2.mem[31][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__B2 (.I(\u2.mem[31][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__I1 (.I(\u2.mem[31][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07895__B2 (.I(\u2.mem[31][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__I1 (.I(\u2.mem[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__B2 (.I(\u2.mem[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__I1 (.I(\u2.mem[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__B2 (.I(\u2.mem[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__I1 (.I(\u2.mem[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__B2 (.I(\u2.mem[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__I1 (.I(\u2.mem[31][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__B2 (.I(\u2.mem[31][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__I1 (.I(\u2.mem[31][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07674__B2 (.I(\u2.mem[31][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__I1 (.I(\u2.mem[32][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07693__A1 (.I(\u2.mem[32][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__I1 (.I(\u2.mem[32][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__A1 (.I(\u2.mem[32][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__I1 (.I(\u2.mem[32][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__A1 (.I(\u2.mem[32][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__I1 (.I(\u2.mem[32][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07867__A1 (.I(\u2.mem[32][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__I1 (.I(\u2.mem[32][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07910__A1 (.I(\u2.mem[32][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__I1 (.I(\u2.mem[32][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07158__A1 (.I(\u2.mem[32][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09500__I1 (.I(\u2.mem[32][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__A1 (.I(\u2.mem[32][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__I1 (.I(\u2.mem[32][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__A1 (.I(\u2.mem[32][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__I1 (.I(\u2.mem[32][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07395__A1 (.I(\u2.mem[32][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__I1 (.I(\u2.mem[32][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__A1 (.I(\u2.mem[32][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__I1 (.I(\u2.mem[32][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07499__A1 (.I(\u2.mem[32][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__I1 (.I(\u2.mem[32][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__A1 (.I(\u2.mem[32][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__I1 (.I(\u2.mem[32][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__A1 (.I(\u2.mem[32][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__I1 (.I(\u2.mem[33][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__B2 (.I(\u2.mem[33][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__I1 (.I(\u2.mem[33][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07562__B2 (.I(\u2.mem[33][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09586__I1 (.I(\u2.mem[34][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06970__B2 (.I(\u2.mem[34][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__I1 (.I(\u2.mem[34][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__B2 (.I(\u2.mem[34][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__I1 (.I(\u2.mem[36][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07022__B2 (.I(\u2.mem[36][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__I1 (.I(\u2.mem[36][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__B2 (.I(\u2.mem[36][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__I1 (.I(\u2.mem[36][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__B2 (.I(\u2.mem[36][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__I1 (.I(\u2.mem[36][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07879__B2 (.I(\u2.mem[36][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__I1 (.I(\u2.mem[36][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__B2 (.I(\u2.mem[36][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__I1 (.I(\u2.mem[36][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07174__B2 (.I(\u2.mem[36][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__I1 (.I(\u2.mem[36][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__B2 (.I(\u2.mem[36][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__I1 (.I(\u2.mem[37][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07064__A1 (.I(\u2.mem[37][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__I1 (.I(\u2.mem[37][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__A1 (.I(\u2.mem[37][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__I1 (.I(\u2.mem[37][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__A1 (.I(\u2.mem[37][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__I1 (.I(\u2.mem[37][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__A1 (.I(\u2.mem[37][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__I1 (.I(\u2.mem[37][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07589__A1 (.I(\u2.mem[37][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__I1 (.I(\u2.mem[38][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07151__B2 (.I(\u2.mem[38][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__I1 (.I(\u2.mem[38][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__B2 (.I(\u2.mem[38][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__I1 (.I(\u2.mem[38][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__B2 (.I(\u2.mem[38][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__I1 (.I(\u2.mem[38][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__B2 (.I(\u2.mem[38][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__I1 (.I(\u2.mem[38][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__B2 (.I(\u2.mem[38][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__I1 (.I(\u2.mem[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07801__A1 (.I(\u2.mem[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__I1 (.I(\u2.mem[40][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A1 (.I(\u2.mem[40][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__I1 (.I(\u2.mem[40][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__A1 (.I(\u2.mem[40][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__I1 (.I(\u2.mem[40][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__A1 (.I(\u2.mem[40][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09886__I1 (.I(\u2.mem[41][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07242__B2 (.I(\u2.mem[41][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__I1 (.I(\u2.mem[41][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07355__B2 (.I(\u2.mem[41][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__I1 (.I(\u2.mem[42][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07470__B2 (.I(\u2.mem[42][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__I1 (.I(\u2.mem[44][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A1 (.I(\u2.mem[44][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__I1 (.I(\u2.mem[45][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07306__A1 (.I(\u2.mem[45][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__I1 (.I(\u2.mem[46][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__B2 (.I(\u2.mem[46][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__I1 (.I(\u2.mem[46][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07883__B2 (.I(\u2.mem[46][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__I1 (.I(\u2.mem[46][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__B2 (.I(\u2.mem[46][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__I1 (.I(\u2.mem[46][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__B2 (.I(\u2.mem[46][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__I1 (.I(\u2.mem[47][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07731__B2 (.I(\u2.mem[47][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__I1 (.I(\u2.mem[47][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__B2 (.I(\u2.mem[47][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__I1 (.I(\u2.mem[48][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07449__B2 (.I(\u2.mem[48][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__I1 (.I(\u2.mem[49][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07814__A1 (.I(\u2.mem[49][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__I1 (.I(\u2.mem[49][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A1 (.I(\u2.mem[49][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__I1 (.I(\u2.mem[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__B2 (.I(\u2.mem[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__I1 (.I(\u2.mem[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__B2 (.I(\u2.mem[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__I1 (.I(\u2.mem[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07859__B2 (.I(\u2.mem[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__I1 (.I(\u2.mem[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__B2 (.I(\u2.mem[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__I1 (.I(\u2.mem[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__B2 (.I(\u2.mem[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08273__I1 (.I(\u2.mem[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__B2 (.I(\u2.mem[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__I1 (.I(\u2.mem[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__B2 (.I(\u2.mem[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__I1 (.I(\u2.mem[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07450__B2 (.I(\u2.mem[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__I1 (.I(\u2.mem[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07622__B2 (.I(\u2.mem[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__I1 (.I(\u2.mem[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__B2 (.I(\u2.mem[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__I1 (.I(\u2.mem[52][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07125__A1 (.I(\u2.mem[52][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__I1 (.I(\u2.mem[52][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__A1 (.I(\u2.mem[52][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__I1 (.I(\u2.mem[52][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__A1 (.I(\u2.mem[52][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__I1 (.I(\u2.mem[52][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07295__A1 (.I(\u2.mem[52][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__I1 (.I(\u2.mem[53][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__A1 (.I(\u2.mem[53][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__I1 (.I(\u2.mem[53][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__A1 (.I(\u2.mem[53][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10428__I1 (.I(\u2.mem[53][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__A1 (.I(\u2.mem[53][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__I1 (.I(\u2.mem[53][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07964__A1 (.I(\u2.mem[53][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__I1 (.I(\u2.mem[53][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__A1 (.I(\u2.mem[53][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__I1 (.I(\u2.mem[53][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__A1 (.I(\u2.mem[53][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__I1 (.I(\u2.mem[53][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__A1 (.I(\u2.mem[53][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__I1 (.I(\u2.mem[53][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__A1 (.I(\u2.mem[53][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__I1 (.I(\u2.mem[55][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__B2 (.I(\u2.mem[55][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10541__I1 (.I(\u2.mem[56][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__B2 (.I(\u2.mem[56][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__I1 (.I(\u2.mem[56][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__B2 (.I(\u2.mem[56][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__I1 (.I(\u2.mem[56][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__B2 (.I(\u2.mem[56][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__I1 (.I(\u2.mem[56][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__B2 (.I(\u2.mem[56][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__I1 (.I(\u2.mem[56][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__B2 (.I(\u2.mem[56][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__I1 (.I(\u2.mem[57][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__A1 (.I(\u2.mem[57][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__I1 (.I(\u2.mem[58][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__A1 (.I(\u2.mem[58][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__I1 (.I(\u2.mem[58][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__A1 (.I(\u2.mem[58][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10609__I1 (.I(\u2.mem[58][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07336__A1 (.I(\u2.mem[58][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__I1 (.I(\u2.mem[58][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__A1 (.I(\u2.mem[58][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__I1 (.I(\u2.mem[58][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07468__A1 (.I(\u2.mem[58][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__I1 (.I(\u2.mem[58][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__A1 (.I(\u2.mem[58][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10620__I1 (.I(\u2.mem[58][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07648__A1 (.I(\u2.mem[58][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__I1 (.I(\u2.mem[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__A1 (.I(\u2.mem[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__I1 (.I(\u2.mem[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__A1 (.I(\u2.mem[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__I1 (.I(\u2.mem[61][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07083__A1 (.I(\u2.mem[61][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__I1 (.I(\u2.mem[61][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__A1 (.I(\u2.mem[61][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__I1 (.I(\u2.mem[61][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__A1 (.I(\u2.mem[61][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__I1 (.I(\u2.mem[61][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07346__A1 (.I(\u2.mem[61][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10729__I1 (.I(\u2.mem[61][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__A1 (.I(\u2.mem[61][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10732__I1 (.I(\u2.mem[61][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__A1 (.I(\u2.mem[61][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10794__I1 (.I(\u2.mem[62][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__B2 (.I(\u2.mem[62][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__I1 (.I(\u2.mem[62][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__B2 (.I(\u2.mem[62][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__I1 (.I(\u2.mem[62][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__B2 (.I(\u2.mem[62][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__I1 (.I(\u2.mem[62][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07428__B2 (.I(\u2.mem[62][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10831__I0 (.I(\u2.mem[63][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07887__B2 (.I(\u2.mem[63][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10835__I0 (.I(\u2.mem[63][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__B2 (.I(\u2.mem[63][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__I1 (.I(\u2.mem[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__A1 (.I(\u2.mem[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__I1 (.I(\u2.mem[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07796__B2 (.I(\u2.mem[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08425__I1 (.I(\u2.mem[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07559__B2 (.I(\u2.mem[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__I1 (.I(\u2.mem[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__A1 (.I(\u2.mem[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__I1 (.I(\u2.mem[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__A1 (.I(\u2.mem[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__I1 (.I(\u2.mem[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A1 (.I(\u2.mem[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__I1 (.I(\u2.mem[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07622__A1 (.I(\u2.mem[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__I1 (.I(\u2.mem[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__A1 (.I(\u2.mem[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__I1 (.I(\u2.mem[9][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__A1 (.I(\u2.mem[9][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__I1 (.I(\u2.mem[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__A1 (.I(\u2.mem[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__I1 (.I(\u2.mem[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__A1 (.I(\u2.mem[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08533__I1 (.I(\u2.mem[9][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__A1 (.I(\u2.mem[9][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__I1 (.I(\u2.mem[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07363__A1 (.I(\u2.mem[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__I1 (.I(\u2.mem[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__A1 (.I(\u2.mem[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__I1 (.I(\u2.mem[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__A1 (.I(\u2.mem[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__A1 (.I(\u3.data ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06036__A1 (.I(\u3.data ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12037__D (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12039__D (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12043__D (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12049__D (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12069__D (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12071__D (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12073__D (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12075__D (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12077__D (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12079__D (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12051__D (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12053__D (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12055__D (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12057__D (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12059__D (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12061__D (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12063__D (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12065__D (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12067__D (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12091__D (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12005__D (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12007__D (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12009__D (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12011__D (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12015__D (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12017__D (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12019__D (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12085__D (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12089__D (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12087__D (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12025__D (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12027__D (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12029__D (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12031__D (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12033__D (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12035__D (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13292__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13285__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13281__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13280__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13282__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13343__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13328__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13330__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13341__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13327__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13329__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13333__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13345__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13342__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13339__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13340__CLK (.I(clknet_leaf_4_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13270__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13271__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13267__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13269__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13334__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13346__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13337__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13278__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13273__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13268__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13338__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13569__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13570__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12133__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13537__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12134__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13553__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13554__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13523__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13524__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13568__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13567__CLK (.I(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13522__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13521__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13563__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13519__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13520__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13565__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13566__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13348__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13336__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13347__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13335__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13574__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13573__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13572__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13571__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13107__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13108__CLK (.I(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13123__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13139__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13542__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13541__CLK (.I(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13140__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13091__CLK (.I(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13124__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13094__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13125__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13126__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13142__CLK (.I(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13076__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13093__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13092__CLK (.I(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13046__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13045__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13075__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13077__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13078__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13061__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12787__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13043__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13044__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13060__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13059__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12710__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12709__CLK (.I(clknet_leaf_27_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13014__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11998__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11999__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12000__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12070__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12072__CLK (.I(clknet_leaf_28_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12950__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12707__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13062__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13029__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12982__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13028__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12981__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12934__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13012__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13576__CLK (.I(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13560__CLK (.I(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13561__CLK (.I(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13543__CLK (.I(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13544__CLK (.I(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12066__CLK (.I(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13030__CLK (.I(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12068__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11997__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12996__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13559__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13575__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13538__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12132__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13540__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13539__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13547__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12129__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12130__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13577__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12131__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12127__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13431__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13378__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12124__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13578__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12136__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12135__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12123__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12128__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13111__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13146__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13546__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12138__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12137__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13143__CLK (.I(clknet_leaf_39_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13144__CLK (.I(clknet_leaf_39_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13145__CLK (.I(clknet_leaf_39_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13112__CLK (.I(clknet_leaf_39_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13562__CLK (.I(clknet_leaf_40_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12004__CLK (.I(clknet_leaf_40_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13081__CLK (.I(clknet_leaf_40_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12979__CLK (.I(clknet_leaf_42_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13027__CLK (.I(clknet_leaf_42_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13082__CLK (.I(clknet_leaf_42_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12001__CLK (.I(clknet_leaf_42_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12002__CLK (.I(clknet_leaf_42_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13079__CLK (.I(clknet_leaf_43_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13080__CLK (.I(clknet_leaf_43_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12730__CLK (.I(clknet_leaf_43_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12727__CLK (.I(clknet_leaf_43_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12980__CLK (.I(clknet_leaf_43_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13050__CLK (.I(clknet_leaf_44_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13048__CLK (.I(clknet_leaf_44_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12792__CLK (.I(clknet_leaf_44_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12791__CLK (.I(clknet_leaf_44_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12729__CLK (.I(clknet_leaf_44_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13047__CLK (.I(clknet_leaf_44_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12951__CLK (.I(clknet_leaf_49_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12714__CLK (.I(clknet_leaf_49_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12935__CLK (.I(clknet_leaf_49_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12952__CLK (.I(clknet_leaf_49_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12746__CLK (.I(clknet_leaf_50_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12713__CLK (.I(clknet_leaf_50_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12712__CLK (.I(clknet_leaf_50_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12744__CLK (.I(clknet_leaf_50_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12759__CLK (.I(clknet_leaf_50_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12218__CLK (.I(clknet_leaf_52_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12231__CLK (.I(clknet_leaf_52_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12234__CLK (.I(clknet_leaf_52_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12215__CLK (.I(clknet_leaf_53_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12217__CLK (.I(clknet_leaf_53_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12743__CLK (.I(clknet_leaf_53_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12745__CLK (.I(clknet_leaf_53_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12202__CLK (.I(clknet_leaf_54_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12201__CLK (.I(clknet_leaf_54_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12728__CLK (.I(clknet_leaf_54_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12265__CLK (.I(clknet_leaf_54_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12248__CLK (.I(clknet_leaf_55_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12249__CLK (.I(clknet_leaf_55_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12266__CLK (.I(clknet_leaf_55_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12263__CLK (.I(clknet_leaf_55_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12247__CLK (.I(clknet_leaf_55_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12666__CLK (.I(clknet_leaf_56_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12154__CLK (.I(clknet_leaf_56_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12153__CLK (.I(clknet_leaf_56_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12888__CLK (.I(clknet_leaf_57_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12887__CLK (.I(clknet_leaf_57_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12250__CLK (.I(clknet_leaf_57_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12233__CLK (.I(clknet_leaf_57_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12232__CLK (.I(clknet_leaf_57_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12665__CLK (.I(clknet_leaf_58_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12663__CLK (.I(clknet_leaf_58_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12106__CLK (.I(clknet_leaf_58_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12375__CLK (.I(clknet_leaf_59_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12346__CLK (.I(clknet_leaf_59_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12184__CLK (.I(clknet_leaf_59_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12185__CLK (.I(clknet_leaf_59_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12186__CLK (.I(clknet_leaf_59_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12819__CLK (.I(clknet_leaf_60_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12916__CLK (.I(clknet_leaf_60_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12867__CLK (.I(clknet_leaf_60_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12377__CLK (.I(clknet_leaf_60_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12345__CLK (.I(clknet_leaf_60_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12378__CLK (.I(clknet_leaf_60_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12836__CLK (.I(clknet_leaf_61_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12183__CLK (.I(clknet_leaf_61_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12820__CLK (.I(clknet_leaf_61_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12884__CLK (.I(clknet_leaf_63_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12886__CLK (.I(clknet_leaf_63_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12885__CLK (.I(clknet_leaf_63_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12104__CLK (.I(clknet_leaf_63_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12105__CLK (.I(clknet_leaf_63_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12838__CLK (.I(clknet_leaf_63_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12227__CLK (.I(clknet_leaf_64_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12152__CLK (.I(clknet_leaf_64_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12151__CLK (.I(clknet_leaf_64_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12883__CLK (.I(clknet_leaf_64_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12899__CLK (.I(clknet_leaf_64_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12755__CLK (.I(clknet_leaf_64_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12228__CLK (.I(clknet_leaf_64_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12740__CLK (.I(clknet_leaf_67_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12949__CLK (.I(clknet_leaf_67_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12212__CLK (.I(clknet_leaf_67_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12933__CLK (.I(clknet_leaf_67_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12213__CLK (.I(clknet_leaf_68_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12214__CLK (.I(clknet_leaf_68_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12708__CLK (.I(clknet_leaf_68_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12756__CLK (.I(clknet_leaf_69_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12262__CLK (.I(clknet_leaf_69_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12230__CLK (.I(clknet_leaf_69_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12229__CLK (.I(clknet_leaf_69_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12742__CLK (.I(clknet_leaf_70_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12741__CLK (.I(clknet_leaf_70_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12261__CLK (.I(clknet_leaf_70_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12259__CLK (.I(clknet_leaf_70_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12260__CLK (.I(clknet_leaf_70_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12757__CLK (.I(clknet_leaf_70_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12723__CLK (.I(clknet_leaf_71_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12790__CLK (.I(clknet_leaf_71_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12789__CLK (.I(clknet_leaf_71_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12196__CLK (.I(clknet_leaf_71_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12788__CLK (.I(clknet_leaf_71_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12195__CLK (.I(clknet_leaf_72_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12197__CLK (.I(clknet_leaf_72_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12724__CLK (.I(clknet_leaf_72_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12725__CLK (.I(clknet_leaf_72_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12726__CLK (.I(clknet_leaf_72_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12147__CLK (.I(clknet_leaf_73_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12150__CLK (.I(clknet_leaf_73_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12149__CLK (.I(clknet_leaf_73_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12246__CLK (.I(clknet_leaf_73_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12243__CLK (.I(clknet_leaf_73_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12198__CLK (.I(clknet_leaf_73_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12245__CLK (.I(clknet_leaf_73_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12902__CLK (.I(clknet_leaf_74_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12901__CLK (.I(clknet_leaf_74_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12758__CLK (.I(clknet_leaf_74_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12244__CLK (.I(clknet_leaf_74_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12148__CLK (.I(clknet_leaf_74_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12660__CLK (.I(clknet_leaf_75_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12180__CLK (.I(clknet_leaf_75_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12900__CLK (.I(clknet_leaf_75_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12661__CLK (.I(clknet_leaf_77_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12339__CLK (.I(clknet_leaf_77_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12387__CLK (.I(clknet_leaf_77_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12390__CLK (.I(clknet_leaf_77_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12182__CLK (.I(clknet_leaf_77_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12181__CLK (.I(clknet_leaf_77_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12342__CLK (.I(clknet_leaf_78_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12374__CLK (.I(clknet_leaf_78_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12371__CLK (.I(clknet_leaf_78_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12389__CLK (.I(clknet_leaf_78_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12358__CLK (.I(clknet_leaf_80_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12356__CLK (.I(clknet_leaf_80_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12357__CLK (.I(clknet_leaf_80_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12869__CLK (.I(clknet_leaf_80_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12853__CLK (.I(clknet_leaf_80_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12854__CLK (.I(clknet_leaf_80_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12372__CLK (.I(clknet_leaf_80_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12340__CLK (.I(clknet_leaf_80_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12917__CLK (.I(clknet_leaf_83_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12868__CLK (.I(clknet_leaf_83_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12870__CLK (.I(clknet_leaf_83_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12355__CLK (.I(clknet_leaf_83_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12821__CLK (.I(clknet_leaf_83_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12822__CLK (.I(clknet_leaf_83_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12452__CLK (.I(clknet_leaf_84_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12324__CLK (.I(clknet_leaf_84_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12451__CLK (.I(clknet_leaf_84_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12323__CLK (.I(clknet_leaf_84_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12918__CLK (.I(clknet_leaf_84_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12454__CLK (.I(clknet_leaf_85_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12326__CLK (.I(clknet_leaf_85_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12325__CLK (.I(clknet_leaf_85_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12965__CLK (.I(clknet_leaf_85_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12677__CLK (.I(clknet_leaf_90_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12771__CLK (.I(clknet_leaf_90_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12852__CLK (.I(clknet_leaf_90_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12676__CLK (.I(clknet_leaf_90_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12164__CLK (.I(clknet_leaf_91_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12165__CLK (.I(clknet_leaf_91_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12166__CLK (.I(clknet_leaf_91_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12163__CLK (.I(clknet_leaf_91_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12772__CLK (.I(clknet_leaf_91_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12518__CLK (.I(clknet_leaf_94_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12563__CLK (.I(clknet_leaf_94_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12643__CLK (.I(clknet_leaf_94_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12613__CLK (.I(clknet_leaf_94_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12611__CLK (.I(clknet_leaf_94_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12566__CLK (.I(clknet_leaf_94_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12565__CLK (.I(clknet_leaf_96_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12630__CLK (.I(clknet_leaf_96_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12598__CLK (.I(clknet_leaf_96_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12534__CLK (.I(clknet_leaf_97_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12629__CLK (.I(clknet_leaf_97_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12627__CLK (.I(clknet_leaf_97_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12628__CLK (.I(clknet_leaf_97_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12581__CLK (.I(clknet_leaf_98_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12580__CLK (.I(clknet_leaf_98_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12532__CLK (.I(clknet_leaf_98_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12550__CLK (.I(clknet_leaf_98_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12548__CLK (.I(clknet_leaf_98_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12549__CLK (.I(clknet_leaf_98_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12533__CLK (.I(clknet_leaf_98_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12582__CLK (.I(clknet_leaf_100_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12308__CLK (.I(clknet_leaf_100_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12309__CLK (.I(clknet_leaf_100_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12485__CLK (.I(clknet_leaf_100_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12486__CLK (.I(clknet_leaf_100_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12278__CLK (.I(clknet_leaf_101_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12292__CLK (.I(clknet_leaf_101_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12294__CLK (.I(clknet_leaf_101_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12293__CLK (.I(clknet_leaf_101_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12275__CLK (.I(clknet_leaf_102_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12276__CLK (.I(clknet_leaf_102_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12277__CLK (.I(clknet_leaf_102_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12531__CLK (.I(clknet_leaf_103_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12633__CLK (.I(clknet_leaf_103_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12547__CLK (.I(clknet_leaf_103_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12291__CLK (.I(clknet_leaf_103_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12632__CLK (.I(clknet_leaf_104_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12307__CLK (.I(clknet_leaf_104_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12579__CLK (.I(clknet_leaf_104_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12595__CLK (.I(clknet_leaf_105_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12484__CLK (.I(clknet_leaf_105_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12468__CLK (.I(clknet_leaf_105_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12515__CLK (.I(clknet_leaf_105_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12500__CLK (.I(clknet_leaf_105_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12470__CLK (.I(clknet_leaf_106_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12469__CLK (.I(clknet_leaf_106_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12502__CLK (.I(clknet_leaf_106_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12501__CLK (.I(clknet_leaf_106_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12420__CLK (.I(clknet_leaf_108_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12435__CLK (.I(clknet_leaf_108_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12403__CLK (.I(clknet_leaf_108_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12467__CLK (.I(clknet_leaf_108_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12170__CLK (.I(clknet_leaf_109_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12167__CLK (.I(clknet_leaf_109_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12168__CLK (.I(clknet_leaf_109_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12963__CLK (.I(clknet_leaf_109_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12964__CLK (.I(clknet_leaf_109_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12650__CLK (.I(clknet_leaf_110_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12419__CLK (.I(clknet_leaf_110_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12698__CLK (.I(clknet_leaf_110_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12695__CLK (.I(clknet_leaf_110_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12618__CLK (.I(clknet_leaf_111_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12697__CLK (.I(clknet_leaf_111_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12570__CLK (.I(clknet_leaf_111_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12617__CLK (.I(clknet_leaf_111_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12649__CLK (.I(clknet_leaf_111_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12522__CLK (.I(clknet_leaf_112_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12407__CLK (.I(clknet_leaf_112_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12410__CLK (.I(clknet_leaf_112_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12568__CLK (.I(clknet_leaf_112_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12426__CLK (.I(clknet_leaf_112_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12616__CLK (.I(clknet_leaf_113_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12615__CLK (.I(clknet_leaf_113_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12599__CLK (.I(clknet_leaf_113_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12602__CLK (.I(clknet_leaf_113_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12567__CLK (.I(clknet_leaf_113_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12569__CLK (.I(clknet_leaf_113_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12634__CLK (.I(clknet_leaf_114_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12631__CLK (.I(clknet_leaf_114_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12648__CLK (.I(clknet_leaf_114_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12647__CLK (.I(clknet_leaf_114_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12538__CLK (.I(clknet_leaf_115_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12535__CLK (.I(clknet_leaf_115_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12551__CLK (.I(clknet_leaf_115_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12583__CLK (.I(clknet_leaf_115_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12586__CLK (.I(clknet_leaf_115_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12584__CLK (.I(clknet_leaf_115_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12585__CLK (.I(clknet_leaf_115_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12601__CLK (.I(clknet_leaf_116_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12536__CLK (.I(clknet_leaf_116_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12537__CLK (.I(clknet_leaf_116_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12313__CLK (.I(clknet_leaf_118_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12314__CLK (.I(clknet_leaf_118_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12311__CLK (.I(clknet_leaf_118_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12520__CLK (.I(clknet_leaf_118_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12521__CLK (.I(clknet_leaf_118_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12282__CLK (.I(clknet_leaf_119_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12281__CLK (.I(clknet_leaf_119_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12554__CLK (.I(clknet_leaf_119_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12552__CLK (.I(clknet_leaf_119_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12553__CLK (.I(clknet_leaf_119_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12295__CLK (.I(clknet_leaf_120_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12296__CLK (.I(clknet_leaf_120_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12280__CLK (.I(clknet_leaf_120_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12297__CLK (.I(clknet_leaf_120_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12279__CLK (.I(clknet_leaf_120_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12472__CLK (.I(clknet_leaf_121_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12490__CLK (.I(clknet_leaf_121_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12506__CLK (.I(clknet_leaf_121_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12489__CLK (.I(clknet_leaf_121_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12503__CLK (.I(clknet_leaf_121_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12312__CLK (.I(clknet_leaf_121_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12487__CLK (.I(clknet_leaf_121_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12504__CLK (.I(clknet_leaf_121_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12499__CLK (.I(clknet_leaf_123_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12483__CLK (.I(clknet_leaf_123_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12474__CLK (.I(clknet_leaf_123_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12424__CLK (.I(clknet_leaf_123_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12440__CLK (.I(clknet_leaf_123_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12968__CLK (.I(clknet_leaf_124_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12970__CLK (.I(clknet_leaf_124_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12434__CLK (.I(clknet_leaf_124_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12967__CLK (.I(clknet_leaf_124_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12919__CLK (.I(clknet_leaf_125_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12329__CLK (.I(clknet_leaf_125_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12969__CLK (.I(clknet_leaf_125_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12330__CLK (.I(clknet_leaf_125_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12457__CLK (.I(clknet_leaf_126_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12456__CLK (.I(clknet_leaf_126_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12328__CLK (.I(clknet_leaf_126_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12327__CLK (.I(clknet_leaf_126_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12922__CLK (.I(clknet_leaf_126_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12441__CLK (.I(clknet_leaf_127_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12458__CLK (.I(clknet_leaf_127_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12439__CLK (.I(clknet_leaf_127_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12682__CLK (.I(clknet_leaf_127_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12455__CLK (.I(clknet_leaf_127_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12442__CLK (.I(clknet_leaf_128_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12423__CLK (.I(clknet_leaf_128_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12425__CLK (.I(clknet_leaf_128_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12856__CLK (.I(clknet_leaf_129_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12858__CLK (.I(clknet_leaf_129_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12681__CLK (.I(clknet_leaf_129_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12696__CLK (.I(clknet_leaf_129_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12680__CLK (.I(clknet_leaf_129_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12778__CLK (.I(clknet_leaf_130_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12777__CLK (.I(clknet_leaf_130_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12679__CLK (.I(clknet_leaf_130_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12776__CLK (.I(clknet_leaf_130_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12392__CLK (.I(clknet_leaf_133_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12359__CLK (.I(clknet_leaf_133_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12361__CLK (.I(clknet_leaf_133_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12857__CLK (.I(clknet_leaf_133_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12855__CLK (.I(clknet_leaf_133_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12839__CLK (.I(clknet_leaf_135_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12823__CLK (.I(clknet_leaf_135_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12108__CLK (.I(clknet_leaf_135_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12664__CLK (.I(clknet_leaf_135_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12107__CLK (.I(clknet_leaf_135_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12871__CLK (.I(clknet_leaf_136_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12360__CLK (.I(clknet_leaf_136_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12825__CLK (.I(clknet_leaf_136_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12826__CLK (.I(clknet_leaf_136_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12840__CLK (.I(clknet_leaf_139_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12808__CLK (.I(clknet_leaf_139_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12810__CLK (.I(clknet_leaf_139_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12809__CLK (.I(clknet_leaf_139_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12842__CLK (.I(clknet_leaf_139_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12903__CLK (.I(clknet_leaf_140_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12890__CLK (.I(clknet_leaf_140_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12109__CLK (.I(clknet_leaf_140_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12807__CLK (.I(clknet_leaf_140_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12761__CLK (.I(clknet_leaf_141_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12905__CLK (.I(clknet_leaf_141_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12906__CLK (.I(clknet_leaf_141_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12881__CLK (.I(clknet_leaf_143_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12226__CLK (.I(clknet_leaf_143_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12803__CLK (.I(clknet_leaf_145_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12802__CLK (.I(clknet_leaf_145_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12834__CLK (.I(clknet_leaf_145_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12832__CLK (.I(clknet_leaf_145_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12818__CLK (.I(clknet_leaf_147_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12912__CLK (.I(clknet_leaf_147_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12816__CLK (.I(clknet_leaf_147_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12915__CLK (.I(clknet_leaf_147_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12351__CLK (.I(clknet_leaf_148_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12833__CLK (.I(clknet_leaf_148_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12352__CLK (.I(clknet_leaf_148_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12863__CLK (.I(clknet_leaf_148_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12864__CLK (.I(clknet_leaf_148_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12865__CLK (.I(clknet_leaf_148_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12850__CLK (.I(clknet_leaf_150_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12354__CLK (.I(clknet_leaf_150_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12370__CLK (.I(clknet_leaf_150_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12353__CLK (.I(clknet_leaf_150_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12848__CLK (.I(clknet_leaf_151_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12847__CLK (.I(clknet_leaf_151_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12866__CLK (.I(clknet_leaf_151_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12337__CLK (.I(clknet_leaf_152_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12160__CLK (.I(clknet_leaf_152_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12335__CLK (.I(clknet_leaf_152_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12338__CLK (.I(clknet_leaf_152_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12769__CLK (.I(clknet_leaf_154_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12849__CLK (.I(clknet_leaf_154_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12674__CLK (.I(clknet_leaf_154_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12673__CLK (.I(clknet_leaf_154_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12161__CLK (.I(clknet_leaf_154_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12402__CLK (.I(clknet_leaf_155_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12959__CLK (.I(clknet_leaf_155_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12399__CLK (.I(clknet_leaf_155_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12609__CLK (.I(clknet_leaf_155_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12768__CLK (.I(clknet_leaf_155_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12767__CLK (.I(clknet_leaf_155_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12770__CLK (.I(clknet_leaf_155_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12961__CLK (.I(clknet_leaf_157_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12914__CLK (.I(clknet_leaf_157_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12319__CLK (.I(clknet_leaf_157_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12911__CLK (.I(clknet_leaf_157_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12321__CLK (.I(clknet_leaf_158_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12913__CLK (.I(clknet_leaf_158_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12322__CLK (.I(clknet_leaf_158_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12320__CLK (.I(clknet_leaf_158_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12432__CLK (.I(clknet_leaf_159_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12450__CLK (.I(clknet_leaf_159_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12447__CLK (.I(clknet_leaf_159_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12448__CLK (.I(clknet_leaf_159_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12921__CLK (.I(clknet_leaf_159_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12449__CLK (.I(clknet_leaf_159_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12401__CLK (.I(clknet_leaf_161_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12417__CLK (.I(clknet_leaf_161_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12498__CLK (.I(clknet_leaf_161_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12433__CLK (.I(clknet_leaf_161_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12513__CLK (.I(clknet_leaf_162_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12514__CLK (.I(clknet_leaf_162_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12512__CLK (.I(clknet_leaf_162_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12511__CLK (.I(clknet_leaf_162_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12466__CLK (.I(clknet_leaf_162_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12505__CLK (.I(clknet_leaf_163_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12497__CLK (.I(clknet_leaf_163_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12496__CLK (.I(clknet_leaf_163_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12495__CLK (.I(clknet_leaf_163_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12479__CLK (.I(clknet_leaf_163_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12488__CLK (.I(clknet_leaf_164_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12482__CLK (.I(clknet_leaf_164_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12287__CLK (.I(clknet_leaf_164_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12304__CLK (.I(clknet_leaf_164_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12305__CLK (.I(clknet_leaf_164_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12480__CLK (.I(clknet_leaf_164_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12481__CLK (.I(clknet_leaf_164_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12273__CLK (.I(clknet_leaf_165_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12288__CLK (.I(clknet_leaf_165_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12290__CLK (.I(clknet_leaf_165_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12298__CLK (.I(clknet_leaf_165_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12289__CLK (.I(clknet_leaf_165_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12303__CLK (.I(clknet_leaf_166_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12306__CLK (.I(clknet_leaf_166_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12271__CLK (.I(clknet_leaf_166_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12529__CLK (.I(clknet_leaf_166_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12530__CLK (.I(clknet_leaf_166_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12274__CLK (.I(clknet_leaf_166_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12272__CLK (.I(clknet_leaf_166_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12543__CLK (.I(clknet_leaf_168_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12544__CLK (.I(clknet_leaf_168_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12545__CLK (.I(clknet_leaf_168_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12546__CLK (.I(clknet_leaf_168_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12592__CLK (.I(clknet_leaf_168_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12624__CLK (.I(clknet_leaf_168_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12559__CLK (.I(clknet_leaf_170_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12561__CLK (.I(clknet_leaf_170_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12299__CLK (.I(clknet_leaf_170_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12577__CLK (.I(clknet_leaf_170_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12626__CLK (.I(clknet_leaf_170_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12463__CLK (.I(clknet_leaf_172_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12608__CLK (.I(clknet_leaf_172_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12640__CLK (.I(clknet_leaf_172_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12623__CLK (.I(clknet_leaf_172_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12591__CLK (.I(clknet_leaf_172_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12625__CLK (.I(clknet_leaf_172_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12641__CLK (.I(clknet_leaf_173_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12607__CLK (.I(clknet_leaf_173_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12610__CLK (.I(clknet_leaf_173_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12464__CLK (.I(clknet_leaf_173_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12398__CLK (.I(clknet_leaf_179_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12510__CLK (.I(clknet_leaf_179_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12507__CLK (.I(clknet_leaf_179_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12459__CLK (.I(clknet_leaf_179_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12395__CLK (.I(clknet_leaf_179_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12509__CLK (.I(clknet_leaf_180_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12508__CLK (.I(clknet_leaf_180_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12396__CLK (.I(clknet_leaf_180_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12397__CLK (.I(clknet_leaf_180_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12428__CLK (.I(clknet_leaf_180_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12478__CLK (.I(clknet_leaf_181_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12494__CLK (.I(clknet_leaf_181_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12302__CLK (.I(clknet_leaf_181_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12300__CLK (.I(clknet_leaf_181_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12477__CLK (.I(clknet_leaf_181_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12476__CLK (.I(clknet_leaf_181_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12571__CLK (.I(clknet_leaf_182_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12491__CLK (.I(clknet_leaf_182_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12475__CLK (.I(clknet_leaf_182_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12575__CLK (.I(clknet_leaf_183_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12523__CLK (.I(clknet_leaf_183_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12301__CLK (.I(clknet_leaf_183_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12284__CLK (.I(clknet_leaf_185_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12285__CLK (.I(clknet_leaf_185_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12286__CLK (.I(clknet_leaf_185_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12268__CLK (.I(clknet_leaf_185_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12270__CLK (.I(clknet_leaf_185_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12269__CLK (.I(clknet_leaf_185_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12524__CLK (.I(clknet_leaf_187_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12526__CLK (.I(clknet_leaf_187_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12573__CLK (.I(clknet_leaf_187_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12589__CLK (.I(clknet_leaf_187_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12541__CLK (.I(clknet_leaf_188_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12525__CLK (.I(clknet_leaf_188_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12542__CLK (.I(clknet_leaf_188_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12622__CLK (.I(clknet_leaf_189_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12540__CLK (.I(clknet_leaf_189_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12492__CLK (.I(clknet_leaf_190_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12590__CLK (.I(clknet_leaf_190_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12588__CLK (.I(clknet_leaf_190_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12621__CLK (.I(clknet_leaf_190_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12620__CLK (.I(clknet_leaf_190_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12556__CLK (.I(clknet_leaf_190_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12638__CLK (.I(clknet_leaf_192_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12636__CLK (.I(clknet_leaf_192_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12557__CLK (.I(clknet_leaf_192_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12637__CLK (.I(clknet_leaf_192_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12669__CLK (.I(clknet_leaf_193_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12668__CLK (.I(clknet_leaf_193_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12684__CLK (.I(clknet_leaf_193_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12685__CLK (.I(clknet_leaf_193_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12686__CLK (.I(clknet_leaf_193_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12606__CLK (.I(clknet_leaf_195_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12683__CLK (.I(clknet_leaf_195_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12667__CLK (.I(clknet_leaf_195_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12429__CLK (.I(clknet_leaf_196_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12460__CLK (.I(clknet_leaf_196_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12957__CLK (.I(clknet_leaf_196_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12603__CLK (.I(clknet_leaf_196_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12461__CLK (.I(clknet_leaf_196_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12605__CLK (.I(clknet_leaf_196_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12317__CLK (.I(clknet_leaf_197_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12958__CLK (.I(clknet_leaf_197_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12956__CLK (.I(clknet_leaf_197_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12413__CLK (.I(clknet_leaf_197_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12843__CLK (.I(clknet_leaf_198_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12955__CLK (.I(clknet_leaf_198_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12412__CLK (.I(clknet_leaf_198_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12445__CLK (.I(clknet_leaf_198_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12444__CLK (.I(clknet_leaf_198_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12318__CLK (.I(clknet_leaf_199_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12862__CLK (.I(clknet_leaf_199_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12859__CLK (.I(clknet_leaf_199_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12446__CLK (.I(clknet_leaf_199_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12443__CLK (.I(clknet_leaf_199_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12350__CLK (.I(clknet_leaf_201_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12812__CLK (.I(clknet_leaf_201_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12813__CLK (.I(clknet_leaf_201_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12910__CLK (.I(clknet_leaf_202_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12909__CLK (.I(clknet_leaf_202_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12908__CLK (.I(clknet_leaf_202_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12348__CLK (.I(clknet_leaf_202_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12349__CLK (.I(clknet_leaf_202_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12764__CLK (.I(clknet_leaf_203_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12846__CLK (.I(clknet_leaf_203_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12766__CLK (.I(clknet_leaf_203_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12763__CLK (.I(clknet_leaf_203_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12860__CLK (.I(clknet_leaf_203_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12653__CLK (.I(clknet_leaf_205_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12654__CLK (.I(clknet_leaf_205_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12380__CLK (.I(clknet_leaf_205_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12158__CLK (.I(clknet_leaf_205_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12652__CLK (.I(clknet_leaf_205_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12157__CLK (.I(clknet_leaf_205_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12845__CLK (.I(clknet_leaf_205_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12156__CLK (.I(clknet_leaf_205_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12334__CLK (.I(clknet_leaf_206_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12332__CLK (.I(clknet_leaf_206_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12364__CLK (.I(clknet_leaf_206_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12381__CLK (.I(clknet_leaf_206_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12829__CLK (.I(clknet_leaf_207_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12331__CLK (.I(clknet_leaf_207_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12379__CLK (.I(clknet_leaf_207_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12651__CLK (.I(clknet_leaf_207_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12382__CLK (.I(clknet_leaf_207_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12333__CLK (.I(clknet_leaf_209_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12366__CLK (.I(clknet_leaf_209_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12892__CLK (.I(clknet_leaf_209_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12171__CLK (.I(clknet_leaf_209_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12174__CLK (.I(clknet_leaf_210_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12173__CLK (.I(clknet_leaf_210_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12172__CLK (.I(clknet_leaf_210_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12365__CLK (.I(clknet_leaf_210_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12748__CLK (.I(clknet_leaf_211_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12235__CLK (.I(clknet_leaf_211_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12204__CLK (.I(clknet_leaf_211_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12238__CLK (.I(clknet_leaf_211_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12237__CLK (.I(clknet_leaf_211_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12236__CLK (.I(clknet_leaf_211_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12140__CLK (.I(clknet_leaf_211_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12141__CLK (.I(clknet_leaf_211_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12142__CLK (.I(clknet_leaf_211_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12206__CLK (.I(clknet_leaf_212_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12205__CLK (.I(clknet_leaf_212_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12749__CLK (.I(clknet_leaf_212_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12139__CLK (.I(clknet_leaf_212_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12750__CLK (.I(clknet_leaf_213_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12221__CLK (.I(clknet_leaf_213_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12253__CLK (.I(clknet_leaf_213_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12877__CLK (.I(clknet_leaf_214_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12894__CLK (.I(clknet_leaf_214_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12095__CLK (.I(clknet_leaf_214_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12096__CLK (.I(clknet_leaf_214_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12893__CLK (.I(clknet_leaf_214_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12252__CLK (.I(clknet_leaf_215_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12220__CLK (.I(clknet_leaf_215_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12876__CLK (.I(clknet_leaf_215_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12731__CLK (.I(clknet_leaf_216_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12251__CLK (.I(clknet_leaf_216_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12747__CLK (.I(clknet_leaf_216_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12222__CLK (.I(clknet_leaf_216_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12254__CLK (.I(clknet_leaf_216_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12219__CLK (.I(clknet_leaf_217_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12239__CLK (.I(clknet_leaf_217_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12203__CLK (.I(clknet_leaf_217_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12255__CLK (.I(clknet_leaf_217_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12094__CLK (.I(clknet_leaf_218_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12177__CLK (.I(clknet_leaf_218_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12175__CLK (.I(clknet_leaf_218_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12143__CLK (.I(clknet_leaf_218_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12145__CLK (.I(clknet_leaf_218_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12875__CLK (.I(clknet_leaf_218_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12795__CLK (.I(clknet_leaf_220_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12814__CLK (.I(clknet_leaf_220_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12830__CLK (.I(clknet_leaf_220_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12798__CLK (.I(clknet_leaf_220_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12797__CLK (.I(clknet_leaf_220_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12796__CLK (.I(clknet_leaf_220_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12907__CLK (.I(clknet_leaf_221_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12811__CLK (.I(clknet_leaf_221_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12347__CLK (.I(clknet_leaf_221_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12384__CLK (.I(clknet_leaf_221_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12827__CLK (.I(clknet_leaf_221_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12656__CLK (.I(clknet_leaf_221_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12383__CLK (.I(clknet_leaf_223_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12655__CLK (.I(clknet_leaf_223_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12385__CLK (.I(clknet_leaf_223_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12369__CLK (.I(clknet_leaf_223_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12367__CLK (.I(clknet_leaf_223_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12896__CLK (.I(clknet_leaf_224_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12897__CLK (.I(clknet_leaf_224_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12098__CLK (.I(clknet_leaf_224_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12657__CLK (.I(clknet_leaf_224_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12658__CLK (.I(clknet_leaf_224_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12386__CLK (.I(clknet_leaf_224_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12242__CLK (.I(clknet_leaf_226_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12144__CLK (.I(clknet_leaf_226_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12176__CLK (.I(clknet_leaf_226_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12241__CLK (.I(clknet_leaf_227_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12240__CLK (.I(clknet_leaf_227_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12752__CLK (.I(clknet_leaf_227_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12193__CLK (.I(clknet_leaf_228_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12256__CLK (.I(clknet_leaf_228_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12258__CLK (.I(clknet_leaf_228_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12257__CLK (.I(clknet_leaf_228_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12192__CLK (.I(clknet_leaf_228_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12882__CLK (.I(clknet_leaf_230_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12880__CLK (.I(clknet_leaf_230_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12879__CLK (.I(clknet_leaf_230_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12898__CLK (.I(clknet_leaf_230_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12753__CLK (.I(clknet_leaf_230_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12208__CLK (.I(clknet_leaf_231_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12223__CLK (.I(clknet_leaf_231_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12224__CLK (.I(clknet_leaf_231_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12931__CLK (.I(clknet_leaf_232_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12225__CLK (.I(clknet_leaf_232_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12210__CLK (.I(clknet_leaf_232_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12209__CLK (.I(clknet_leaf_232_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12737__CLK (.I(clknet_leaf_232_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12929__CLK (.I(clknet_leaf_233_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12945__CLK (.I(clknet_leaf_233_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12946__CLK (.I(clknet_leaf_233_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12947__CLK (.I(clknet_leaf_233_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12721__CLK (.I(clknet_leaf_235_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12722__CLK (.I(clknet_leaf_235_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12928__CLK (.I(clknet_leaf_235_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12785__CLK (.I(clknet_leaf_235_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12944__CLK (.I(clknet_leaf_235_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12994__CLK (.I(clknet_leaf_236_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12720__CLK (.I(clknet_leaf_236_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12719__CLK (.I(clknet_leaf_236_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13073__CLK (.I(clknet_leaf_236_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12191__CLK (.I(clknet_leaf_237_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12735__CLK (.I(clknet_leaf_237_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12943__CLK (.I(clknet_leaf_237_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13010__CLK (.I(clknet_leaf_237_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12704__CLK (.I(clknet_leaf_238_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12706__CLK (.I(clknet_leaf_238_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12705__CLK (.I(clknet_leaf_238_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12194__CLK (.I(clknet_leaf_238_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12991__CLK (.I(clknet_leaf_239_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13009__CLK (.I(clknet_leaf_239_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12993__CLK (.I(clknet_leaf_239_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12703__CLK (.I(clknet_leaf_239_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13071__CLK (.I(clknet_leaf_240_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12992__CLK (.I(clknet_leaf_240_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13008__CLK (.I(clknet_leaf_240_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13057__CLK (.I(clknet_leaf_240_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13007__CLK (.I(clknet_leaf_240_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13055__CLK (.I(clknet_leaf_240_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13106__CLK (.I(clknet_leaf_241_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13089__CLK (.I(clknet_leaf_241_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13072__CLK (.I(clknet_leaf_241_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13074__CLK (.I(clknet_leaf_241_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13058__CLK (.I(clknet_leaf_242_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13090__CLK (.I(clknet_leaf_242_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13122__CLK (.I(clknet_leaf_242_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13104__CLK (.I(clknet_leaf_243_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13119__CLK (.I(clknet_leaf_243_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13056__CLK (.I(clknet_leaf_243_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13088__CLK (.I(clknet_leaf_245_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13087__CLK (.I(clknet_leaf_245_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13099__CLK (.I(clknet_leaf_245_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13152__CLK (.I(clknet_leaf_245_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12987__CLK (.I(clknet_leaf_248_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13067__CLK (.I(clknet_leaf_248_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13035__CLK (.I(clknet_leaf_248_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13038__CLK (.I(clknet_leaf_248_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13023__CLK (.I(clknet_leaf_249_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12975__CLK (.I(clknet_leaf_249_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13019__CLK (.I(clknet_leaf_249_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12976__CLK (.I(clknet_leaf_249_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13003__CLK (.I(clknet_leaf_249_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12939__CLK (.I(clknet_leaf_251_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13025__CLK (.I(clknet_leaf_251_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12187__CLK (.I(clknet_leaf_251_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13026__CLK (.I(clknet_leaf_251_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12715__CLK (.I(clknet_leaf_252_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12718__CLK (.I(clknet_leaf_252_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12734__CLK (.I(clknet_leaf_252_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12189__CLK (.I(clknet_leaf_252_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12188__CLK (.I(clknet_leaf_252_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12190__CLK (.I(clknet_leaf_252_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12923__CLK (.I(clknet_leaf_252_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13070__CLK (.I(clknet_leaf_253_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12780__CLK (.I(clknet_leaf_253_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12781__CLK (.I(clknet_leaf_253_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12782__CLK (.I(clknet_leaf_253_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12779__CLK (.I(clknet_leaf_253_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12717__CLK (.I(clknet_leaf_254_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12716__CLK (.I(clknet_leaf_254_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13051__CLK (.I(clknet_leaf_254_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13068__CLK (.I(clknet_leaf_254_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12700__CLK (.I(clknet_leaf_256_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12940__CLK (.I(clknet_leaf_256_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12702__CLK (.I(clknet_leaf_256_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12941__CLK (.I(clknet_leaf_256_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13004__CLK (.I(clknet_leaf_257_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12988__CLK (.I(clknet_leaf_257_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12925__CLK (.I(clknet_leaf_257_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12924__CLK (.I(clknet_leaf_257_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12701__CLK (.I(clknet_leaf_257_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12990__CLK (.I(clknet_leaf_258_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13020__CLK (.I(clknet_leaf_258_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13021__CLK (.I(clknet_leaf_258_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13005__CLK (.I(clknet_leaf_258_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12989__CLK (.I(clknet_leaf_258_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13053__CLK (.I(clknet_leaf_259_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13069__CLK (.I(clknet_leaf_259_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13054__CLK (.I(clknet_leaf_259_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13052__CLK (.I(clknet_leaf_259_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13006__CLK (.I(clknet_leaf_259_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13022__CLK (.I(clknet_leaf_259_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12974__CLK (.I(clknet_leaf_261_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13084__CLK (.I(clknet_leaf_261_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13155__CLK (.I(clknet_leaf_261_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13116__CLK (.I(clknet_leaf_261_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13117__CLK (.I(clknet_leaf_261_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13168__CLK (.I(clknet_leaf_263_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13173__CLK (.I(clknet_leaf_263_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13172__CLK (.I(clknet_leaf_263_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13167__CLK (.I(clknet_leaf_263_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13166__CLK (.I(clknet_leaf_263_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13154__CLK (.I(clknet_leaf_263_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13148__CLK (.I(clknet_leaf_263_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13171__CLK (.I(clknet_leaf_264_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13165__CLK (.I(clknet_leaf_264_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13100__CLK (.I(clknet_leaf_264_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13149__CLK (.I(clknet_leaf_264_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13132__CLK (.I(clknet_leaf_267_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13083__CLK (.I(clknet_leaf_267_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13086__CLK (.I(clknet_leaf_267_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13037__CLK (.I(clknet_leaf_267_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13170__CLK (.I(clknet_leaf_268_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13153__CLK (.I(clknet_leaf_268_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13133__CLK (.I(clknet_leaf_268_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13134__CLK (.I(clknet_leaf_268_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13188__CLK (.I(clknet_leaf_270_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13164__CLK (.I(clknet_leaf_270_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13264__CLK (.I(clknet_leaf_270_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13261__CLK (.I(clknet_leaf_270_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13262__CLK (.I(clknet_leaf_271_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13206__CLK (.I(clknet_leaf_271_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13200__CLK (.I(clknet_leaf_271_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13181__CLK (.I(clknet_leaf_271_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13182__CLK (.I(clknet_leaf_271_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13246__CLK (.I(clknet_leaf_272_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13241__CLK (.I(clknet_leaf_272_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13235__CLK (.I(clknet_leaf_272_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13194__CLK (.I(clknet_leaf_272_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13263__CLK (.I(clknet_leaf_272_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13248__CLK (.I(clknet_leaf_272_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13247__CLK (.I(clknet_leaf_272_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13159__CLK (.I(clknet_leaf_274_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13163__CLK (.I(clknet_leaf_274_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13187__CLK (.I(clknet_leaf_274_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13193__CLK (.I(clknet_leaf_274_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13199__CLK (.I(clknet_leaf_274_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13179__CLK (.I(clknet_leaf_275_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13174__CLK (.I(clknet_leaf_275_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13180__CLK (.I(clknet_leaf_275_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13162__CLK (.I(clknet_leaf_275_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13205__CLK (.I(clknet_leaf_275_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13177__CLK (.I(clknet_leaf_275_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13186__CLK (.I(clknet_leaf_276_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13204__CLK (.I(clknet_leaf_276_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13198__CLK (.I(clknet_leaf_276_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13192__CLK (.I(clknet_leaf_276_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13160__CLK (.I(clknet_leaf_276_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13178__CLK (.I(clknet_leaf_276_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13161__CLK (.I(clknet_leaf_276_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13190__CLK (.I(clknet_leaf_279_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13191__CLK (.I(clknet_leaf_279_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13232__CLK (.I(clknet_leaf_279_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13230__CLK (.I(clknet_leaf_279_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13227__CLK (.I(clknet_leaf_279_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13226__CLK (.I(clknet_leaf_279_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13222__CLK (.I(clknet_leaf_280_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13228__CLK (.I(clknet_leaf_280_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13202__CLK (.I(clknet_leaf_280_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13203__CLK (.I(clknet_leaf_280_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13221__CLK (.I(clknet_leaf_281_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13208__CLK (.I(clknet_leaf_281_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13210__CLK (.I(clknet_leaf_281_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13209__CLK (.I(clknet_leaf_281_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13225__CLK (.I(clknet_leaf_283_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13218__CLK (.I(clknet_leaf_283_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13219__CLK (.I(clknet_leaf_283_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13215__CLK (.I(clknet_leaf_283_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13249__CLK (.I(clknet_leaf_285_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13250__CLK (.I(clknet_leaf_285_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13251__CLK (.I(clknet_leaf_285_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13233__CLK (.I(clknet_leaf_285_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13245__CLK (.I(clknet_leaf_285_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13217__CLK (.I(clknet_leaf_286_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13224__CLK (.I(clknet_leaf_286_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13229__CLK (.I(clknet_leaf_286_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13223__CLK (.I(clknet_leaf_286_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12052__CLK (.I(clknet_leaf_287_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12054__CLK (.I(clknet_leaf_287_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13211__CLK (.I(clknet_leaf_287_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12022__CLK (.I(clknet_leaf_287_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13207__CLK (.I(clknet_leaf_287_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13480__CLK (.I(clknet_leaf_289_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12034__CLK (.I(clknet_leaf_289_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13485__CLK (.I(clknet_leaf_289_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12024__CLK (.I(clknet_leaf_289_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12020__CLK (.I(clknet_leaf_289_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12014__CLK (.I(clknet_leaf_289_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13479__CLK (.I(clknet_leaf_290_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13478__CLK (.I(clknet_leaf_290_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13484__CLK (.I(clknet_leaf_290_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13483__CLK (.I(clknet_leaf_290_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13254__CLK (.I(clknet_leaf_291_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13252__CLK (.I(clknet_leaf_291_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13212__CLK (.I(clknet_leaf_291_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13243__CLK (.I(clknet_leaf_291_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13253__CLK (.I(clknet_leaf_291_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13244__CLK (.I(clknet_leaf_291_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13492__CLK (.I(clknet_leaf_292_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13490__CLK (.I(clknet_leaf_292_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13491__CLK (.I(clknet_leaf_292_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13473__CLK (.I(clknet_leaf_292_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13494__CLK (.I(clknet_leaf_295_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13476__CLK (.I(clknet_leaf_295_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13475__CLK (.I(clknet_leaf_295_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13260__CLK (.I(clknet_leaf_295_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13266__CLK (.I(clknet_leaf_295_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13265__CLK (.I(clknet_leaf_295_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13255__CLK (.I(clknet_leaf_295_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12088__CLK (.I(clknet_leaf_298_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13420__CLK (.I(clknet_leaf_298_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13486__CLK (.I(clknet_leaf_298_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13477__CLK (.I(clknet_leaf_298_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13488__CLK (.I(clknet_leaf_298_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13482__CLK (.I(clknet_leaf_298_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13417__CLK (.I(clknet_leaf_298_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13402__CLK (.I(clknet_leaf_298_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12042__CLK (.I(clknet_leaf_299_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12040__CLK (.I(clknet_leaf_299_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12018__CLK (.I(clknet_leaf_299_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12044__CLK (.I(clknet_leaf_299_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12008__CLK (.I(clknet_leaf_299_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13418__CLK (.I(clknet_leaf_299_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13316__CLK (.I(clknet_leaf_300_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13315__CLK (.I(clknet_leaf_300_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13454__CLK (.I(clknet_leaf_300_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12058__CLK (.I(clknet_leaf_300_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12064__CLK (.I(clknet_leaf_300_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12060__CLK (.I(clknet_leaf_300_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13453__CLK (.I(clknet_leaf_301_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13317__CLK (.I(clknet_leaf_301_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13319__CLK (.I(clknet_leaf_301_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13383__CLK (.I(clknet_leaf_301_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13384__CLK (.I(clknet_leaf_301_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13318__CLK (.I(clknet_leaf_301_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13400__CLK (.I(clknet_leaf_301_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12032__CLK (.I(clknet_leaf_302_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13455__CLK (.I(clknet_leaf_302_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12092__CLK (.I(clknet_leaf_302_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12062__CLK (.I(clknet_leaf_302_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12038__CLK (.I(clknet_leaf_302_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12026__CLK (.I(clknet_leaf_302_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13323__CLK (.I(clknet_leaf_303_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13321__CLK (.I(clknet_leaf_303_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12080__CLK (.I(clknet_leaf_303_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12090__CLK (.I(clknet_leaf_303_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13457__CLK (.I(clknet_leaf_304_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13405__CLK (.I(clknet_leaf_304_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13456__CLK (.I(clknet_leaf_304_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13326__CLK (.I(clknet_leaf_304_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13408__CLK (.I(clknet_leaf_304_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13407__CLK (.I(clknet_leaf_304_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13406__CLK (.I(clknet_leaf_304_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13409__CLK (.I(clknet_leaf_305_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13404__CLK (.I(clknet_leaf_305_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13381__CLK (.I(clknet_leaf_305_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13410__CLK (.I(clknet_leaf_305_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13458__CLK (.I(clknet_leaf_306_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13385__CLK (.I(clknet_leaf_306_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13386__CLK (.I(clknet_leaf_306_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13320__CLK (.I(clknet_leaf_306_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13395__CLK (.I(clknet_leaf_307_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13397__CLK (.I(clknet_leaf_307_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13398__CLK (.I(clknet_leaf_307_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12028__CLK (.I(clknet_leaf_307_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12030__CLK (.I(clknet_leaf_307_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13256__CLK (.I(clknet_leaf_311_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13259__CLK (.I(clknet_leaf_311_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12036__CLK (.I(clknet_leaf_311_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13103__CLK (.I(clknet_leaf_312_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13496__CLK (.I(clknet_leaf_312_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13258__CLK (.I(clknet_leaf_312_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12006__CLK (.I(clknet_leaf_312_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12010__CLK (.I(clknet_leaf_312_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13257__CLK (.I(clknet_leaf_312_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13138__CLK (.I(clknet_leaf_314_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13121__CLK (.I(clknet_leaf_314_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13105__CLK (.I(clknet_leaf_314_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13135__CLK (.I(clknet_leaf_314_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13526__CLK (.I(clknet_leaf_314_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13529__CLK (.I(clknet_leaf_316_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13527__CLK (.I(clknet_leaf_316_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13497__CLK (.I(clknet_leaf_316_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13499__CLK (.I(clknet_leaf_316_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13530__CLK (.I(clknet_leaf_317_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13511__CLK (.I(clknet_leaf_317_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13500__CLK (.I(clknet_leaf_317_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13528__CLK (.I(clknet_leaf_317_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11989__CLK (.I(clknet_leaf_318_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13534__CLK (.I(clknet_leaf_318_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11991__CLK (.I(clknet_leaf_318_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11993__CLK (.I(clknet_leaf_318_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13536__CLK (.I(clknet_leaf_318_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13517__CLK (.I(clknet_leaf_318_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13533__CLK (.I(clknet_leaf_318_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13505__CLK (.I(clknet_leaf_318_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11995__CLK (.I(clknet_leaf_319_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13017__CLK (.I(clknet_leaf_319_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13016__CLK (.I(clknet_leaf_319_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12985__CLK (.I(clknet_leaf_319_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12784__CLK (.I(clknet_leaf_321_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12786__CLK (.I(clknet_leaf_321_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13041__CLK (.I(clknet_leaf_321_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13042__CLK (.I(clknet_leaf_321_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13000__CLK (.I(clknet_leaf_322_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13018__CLK (.I(clknet_leaf_322_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13001__CLK (.I(clknet_leaf_322_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13002__CLK (.I(clknet_leaf_322_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12783__CLK (.I(clknet_leaf_322_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12937__CLK (.I(clknet_leaf_323_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13011__CLK (.I(clknet_leaf_323_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12995__CLK (.I(clknet_leaf_323_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12999__CLK (.I(clknet_leaf_323_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13015__CLK (.I(clknet_leaf_323_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12954__CLK (.I(clknet_leaf_324_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12936__CLK (.I(clknet_leaf_324_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12953__CLK (.I(clknet_leaf_324_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13034__CLK (.I(clknet_leaf_326_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13031__CLK (.I(clknet_leaf_326_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12986__CLK (.I(clknet_leaf_326_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12983__CLK (.I(clknet_leaf_326_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13129__CLK (.I(clknet_leaf_327_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13113__CLK (.I(clknet_leaf_327_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13127__CLK (.I(clknet_leaf_327_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13130__CLK (.I(clknet_leaf_327_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13032__CLK (.I(clknet_leaf_328_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13033__CLK (.I(clknet_leaf_328_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12122__CLK (.I(clknet_leaf_328_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12116__CLK (.I(clknet_leaf_328_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12121__CLK (.I(clknet_leaf_328_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11990__CLK (.I(clknet_leaf_329_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13535__CLK (.I(clknet_leaf_329_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11992__CLK (.I(clknet_leaf_329_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12984__CLK (.I(clknet_leaf_329_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13501__CLK (.I(clknet_leaf_330_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13507__CLK (.I(clknet_leaf_330_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13506__CLK (.I(clknet_leaf_330_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13512__CLK (.I(clknet_leaf_330_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13518__CLK (.I(clknet_leaf_330_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13504__CLK (.I(clknet_leaf_331_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13508__CLK (.I(clknet_leaf_331_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13502__CLK (.I(clknet_leaf_331_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13503__CLK (.I(clknet_leaf_331_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12113__CLK (.I(clknet_leaf_331_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12115__CLK (.I(clknet_leaf_332_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12119__CLK (.I(clknet_leaf_332_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12111__CLK (.I(clknet_leaf_332_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12117__CLK (.I(clknet_leaf_332_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13433__CLK (.I(clknet_leaf_338_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13516__CLK (.I(clknet_leaf_338_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13411__CLK (.I(clknet_leaf_341_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13416__CLK (.I(clknet_leaf_341_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13439__CLK (.I(clknet_leaf_341_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13440__CLK (.I(clknet_leaf_341_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13322__CLK (.I(clknet_leaf_342_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13324__CLK (.I(clknet_leaf_342_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13451__CLK (.I(clknet_leaf_342_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13414__CLK (.I(clknet_leaf_342_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13452__CLK (.I(clknet_leaf_342_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13325__CLK (.I(clknet_leaf_342_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13415__CLK (.I(clknet_leaf_342_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12076__CLK (.I(clknet_leaf_343_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12078__CLK (.I(clknet_leaf_343_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13448__CLK (.I(clknet_leaf_343_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13447__CLK (.I(clknet_leaf_343_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13449__CLK (.I(clknet_leaf_343_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12074__CLK (.I(clknet_leaf_343_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13450__CLK (.I(clknet_leaf_343_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13464__CLK (.I(clknet_leaf_344_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13413__CLK (.I(clknet_leaf_344_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13412__CLK (.I(clknet_leaf_344_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13463__CLK (.I(clknet_leaf_344_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13461__CLK (.I(clknet_leaf_344_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13467__CLK (.I(clknet_leaf_346_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13465__CLK (.I(clknet_leaf_346_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13468__CLK (.I(clknet_leaf_346_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13462__CLK (.I(clknet_leaf_346_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13311__CLK (.I(clknet_leaf_347_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13466__CLK (.I(clknet_leaf_347_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13424__CLK (.I(clknet_leaf_347_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13470__CLK (.I(clknet_leaf_347_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13423__CLK (.I(clknet_leaf_348_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13441__CLK (.I(clknet_leaf_348_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13309__CLK (.I(clknet_leaf_348_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13312__CLK (.I(clknet_leaf_348_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13310__CLK (.I(clknet_leaf_348_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13427__CLK (.I(clknet_leaf_349_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13426__CLK (.I(clknet_leaf_349_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13314__CLK (.I(clknet_leaf_349_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13444__CLK (.I(clknet_leaf_349_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13313__CLK (.I(clknet_leaf_349_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13425__CLK (.I(clknet_leaf_349_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13445__CLK (.I(clknet_leaf_350_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13436__CLK (.I(clknet_leaf_350_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13446__CLK (.I(clknet_leaf_350_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13435__CLK (.I(clknet_leaf_350_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13437__CLK (.I(clknet_leaf_350_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13428__CLK (.I(clknet_leaf_350_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13362__CLK (.I(clknet_leaf_354_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13373__CLK (.I(clknet_leaf_354_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13367__CLK (.I(clknet_leaf_354_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13290__CLK (.I(clknet_leaf_354_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13387__CLK (.I(clknet_leaf_355_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13390__CLK (.I(clknet_leaf_355_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13388__CLK (.I(clknet_leaf_355_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13361__CLK (.I(clknet_leaf_355_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13389__CLK (.I(clknet_leaf_355_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13374__CLK (.I(clknet_leaf_355_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13358__CLK (.I(clknet_leaf_356_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13369__CLK (.I(clknet_leaf_356_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13442__CLK (.I(clknet_leaf_356_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13443__CLK (.I(clknet_leaf_356_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13357__CLK (.I(clknet_leaf_356_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13360__CLK (.I(clknet_leaf_356_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13359__CLK (.I(clknet_leaf_357_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13371__CLK (.I(clknet_leaf_357_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13370__CLK (.I(clknet_leaf_357_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13353__CLK (.I(clknet_leaf_358_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13305__CLK (.I(clknet_leaf_358_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13306__CLK (.I(clknet_leaf_358_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13365__CLK (.I(clknet_leaf_358_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13364__CLK (.I(clknet_leaf_358_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13363__CLK (.I(clknet_leaf_358_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13307__CLK (.I(clknet_leaf_359_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13368__CLK (.I(clknet_leaf_359_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13372__CLK (.I(clknet_leaf_359_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13366__CLK (.I(clknet_leaf_359_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13354__CLK (.I(clknet_leaf_359_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13283__CLK (.I(clknet_leaf_360_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13355__CLK (.I(clknet_leaf_360_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13356__CLK (.I(clknet_leaf_360_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13351__CLK (.I(clknet_leaf_361_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13352__CLK (.I(clknet_leaf_361_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13291__CLK (.I(clknet_leaf_361_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13279__CLK (.I(clknet_leaf_361_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13299__CLK (.I(clknet_leaf_363_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12093__CLK (.I(clknet_leaf_363_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12083__CLK (.I(clknet_leaf_363_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12084__CLK (.I(clknet_leaf_363_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12082__CLK (.I(clknet_leaf_363_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13297__CLK (.I(clknet_leaf_363_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13288__CLK (.I(clknet_leaf_364_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13294__CLK (.I(clknet_leaf_364_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13287__CLK (.I(clknet_leaf_364_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13293__CLK (.I(clknet_leaf_364_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_1_0_clock_I (.I(clknet_3_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_0_0_clock_I (.I(clknet_3_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_3_0_clock_I (.I(clknet_3_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_2_0_clock_I (.I(clknet_3_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_5_0_clock_I (.I(clknet_3_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_4_0_clock_I (.I(clknet_3_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_7_0_clock_I (.I(clknet_3_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_6_0_clock_I (.I(clknet_3_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_9_0_clock_I (.I(clknet_3_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_8_0_clock_I (.I(clknet_3_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_11_0_clock_I (.I(clknet_3_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_10_0_clock_I (.I(clknet_3_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_13_0_clock_I (.I(clknet_3_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_12_0_clock_I (.I(clknet_3_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_15_0_clock_I (.I(clknet_3_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_14_0_clock_I (.I(clknet_3_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_1_0_clock_I (.I(clknet_4_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_0_0_clock_I (.I(clknet_4_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_3_0_clock_I (.I(clknet_4_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_2_0_clock_I (.I(clknet_4_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_5_0_clock_I (.I(clknet_4_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_4_0_clock_I (.I(clknet_4_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_7_0_clock_I (.I(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_6_0_clock_I (.I(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_9_0_clock_I (.I(clknet_4_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_8_0_clock_I (.I(clknet_4_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_11_0_clock_I (.I(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_10_0_clock_I (.I(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_13_0_clock_I (.I(clknet_4_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_12_0_clock_I (.I(clknet_4_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_15_0_clock_I (.I(clknet_4_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_14_0_clock_I (.I(clknet_4_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_17_0_clock_I (.I(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_16_0_clock_I (.I(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_19_0_clock_I (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_18_0_clock_I (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_21_0_clock_I (.I(clknet_4_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_20_0_clock_I (.I(clknet_4_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_23_0_clock_I (.I(clknet_4_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_22_0_clock_I (.I(clknet_4_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_25_0_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_24_0_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_27_0_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_26_0_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_29_0_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_28_0_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_31_0_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_30_0_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_364_clock_I (.I(clknet_5_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_363_clock_I (.I(clknet_5_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_362_clock_I (.I(clknet_5_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_361_clock_I (.I(clknet_5_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_360_clock_I (.I(clknet_5_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_clock_I (.I(clknet_5_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13272__CLK (.I(clknet_5_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_clock_I (.I(clknet_5_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_clock_I (.I(clknet_5_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_clock_I (.I(clknet_5_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_clock_I (.I(clknet_5_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_clock_I (.I(clknet_5_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_clock_I (.I(clknet_5_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_359_clock_I (.I(clknet_5_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_358_clock_I (.I(clknet_5_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_357_clock_I (.I(clknet_5_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_356_clock_I (.I(clknet_5_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_355_clock_I (.I(clknet_5_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_354_clock_I (.I(clknet_5_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_353_clock_I (.I(clknet_5_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_352_clock_I (.I(clknet_5_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_clock_I (.I(clknet_5_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_clock_I (.I(clknet_5_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_clock_I (.I(clknet_5_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_clock_I (.I(clknet_5_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_clock_I (.I(clknet_5_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_clock_I (.I(clknet_5_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_clock_I (.I(clknet_5_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_clock_I (.I(clknet_5_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_clock_I (.I(clknet_5_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_clock_I (.I(clknet_5_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_clock_I (.I(clknet_5_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_clock_I (.I(clknet_5_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_clock_I (.I(clknet_5_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_clock_I (.I(clknet_5_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_clock_I (.I(clknet_5_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_clock_I (.I(clknet_5_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_clock_I (.I(clknet_5_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_clock_I (.I(clknet_5_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_clock_I (.I(clknet_5_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_clock_I (.I(clknet_5_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_clock_I (.I(clknet_5_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_clock_I (.I(clknet_5_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_clock_I (.I(clknet_5_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_clock_I (.I(clknet_5_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_clock_I (.I(clknet_5_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_clock_I (.I(clknet_5_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_clock_I (.I(clknet_5_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_clock_I (.I(clknet_5_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_clock_I (.I(clknet_5_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13430__CLK (.I(clknet_5_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_350_clock_I (.I(clknet_5_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_349_clock_I (.I(clknet_5_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_348_clock_I (.I(clknet_5_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_347_clock_I (.I(clknet_5_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_346_clock_I (.I(clknet_5_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_337_clock_I (.I(clknet_5_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_336_clock_I (.I(clknet_5_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_clock_I (.I(clknet_5_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_345_clock_I (.I(clknet_5_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_344_clock_I (.I(clknet_5_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_343_clock_I (.I(clknet_5_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_342_clock_I (.I(clknet_5_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_341_clock_I (.I(clknet_5_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_340_clock_I (.I(clknet_5_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13438__CLK (.I(clknet_5_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_338_clock_I (.I(clknet_5_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_335_clock_I (.I(clknet_5_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_334_clock_I (.I(clknet_5_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_333_clock_I (.I(clknet_5_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_clock_I (.I(clknet_5_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_clock_I (.I(clknet_5_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_clock_I (.I(clknet_5_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_clock_I (.I(clknet_5_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_clock_I (.I(clknet_5_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_clock_I (.I(clknet_5_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_clock_I (.I(clknet_5_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_clock_I (.I(clknet_5_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_clock_I (.I(clknet_5_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_332_clock_I (.I(clknet_5_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_331_clock_I (.I(clknet_5_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_330_clock_I (.I(clknet_5_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_329_clock_I (.I(clknet_5_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_328_clock_I (.I(clknet_5_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_327_clock_I (.I(clknet_5_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_326_clock_I (.I(clknet_5_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_325_clock_I (.I(clknet_5_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_324_clock_I (.I(clknet_5_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_clock_I (.I(clknet_5_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_clock_I (.I(clknet_5_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_clock_I (.I(clknet_5_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_clock_I (.I(clknet_5_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_clock_I (.I(clknet_5_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_clock_I (.I(clknet_5_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_clock_I (.I(clknet_5_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_clock_I (.I(clknet_5_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_clock_I (.I(clknet_5_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_clock_I (.I(clknet_5_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_clock_I (.I(clknet_5_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_clock_I (.I(clknet_5_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_clock_I (.I(clknet_5_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_clock_I (.I(clknet_5_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_clock_I (.I(clknet_5_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_clock_I (.I(clknet_5_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_clock_I (.I(clknet_5_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_clock_I (.I(clknet_5_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_clock_I (.I(clknet_5_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_clock_I (.I(clknet_5_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_clock_I (.I(clknet_5_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_clock_I (.I(clknet_5_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_clock_I (.I(clknet_5_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_clock_I (.I(clknet_5_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_clock_I (.I(clknet_5_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_clock_I (.I(clknet_5_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_clock_I (.I(clknet_5_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_clock_I (.I(clknet_5_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_clock_I (.I(clknet_5_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_clock_I (.I(clknet_5_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_clock_I (.I(clknet_5_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_clock_I (.I(clknet_5_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_clock_I (.I(clknet_5_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_clock_I (.I(clknet_5_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_clock_I (.I(clknet_5_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_clock_I (.I(clknet_5_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_clock_I (.I(clknet_5_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_clock_I (.I(clknet_5_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_109_clock_I (.I(clknet_5_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_108_clock_I (.I(clknet_5_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_clock_I (.I(clknet_5_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_clock_I (.I(clknet_5_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_clock_I (.I(clknet_5_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_clock_I (.I(clknet_5_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_clock_I (.I(clknet_5_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_clock_I (.I(clknet_5_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_clock_I (.I(clknet_5_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_clock_I (.I(clknet_5_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_clock_I (.I(clknet_5_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_clock_I (.I(clknet_5_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_clock_I (.I(clknet_5_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_clock_I (.I(clknet_5_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_134_clock_I (.I(clknet_5_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_133_clock_I (.I(clknet_5_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_132_clock_I (.I(clknet_5_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_131_clock_I (.I(clknet_5_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_clock_I (.I(clknet_5_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_clock_I (.I(clknet_5_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_clock_I (.I(clknet_5_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_clock_I (.I(clknet_5_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_clock_I (.I(clknet_5_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_clock_I (.I(clknet_5_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_clock_I (.I(clknet_5_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_clock_I (.I(clknet_5_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_clock_I (.I(clknet_5_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12762__CLK (.I(clknet_5_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_141_clock_I (.I(clknet_5_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_140_clock_I (.I(clknet_5_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_139_clock_I (.I(clknet_5_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_138_clock_I (.I(clknet_5_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_137_clock_I (.I(clknet_5_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_136_clock_I (.I(clknet_5_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_135_clock_I (.I(clknet_5_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_clock_I (.I(clknet_5_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_clock_I (.I(clknet_5_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_130_clock_I (.I(clknet_5_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_129_clock_I (.I(clknet_5_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_128_clock_I (.I(clknet_5_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_117_clock_I (.I(clknet_5_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_116_clock_I (.I(clknet_5_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_115_clock_I (.I(clknet_5_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_114_clock_I (.I(clknet_5_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_113_clock_I (.I(clknet_5_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_112_clock_I (.I(clknet_5_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_111_clock_I (.I(clknet_5_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_110_clock_I (.I(clknet_5_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_127_clock_I (.I(clknet_5_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_126_clock_I (.I(clknet_5_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_125_clock_I (.I(clknet_5_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_124_clock_I (.I(clknet_5_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_123_clock_I (.I(clknet_5_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_122_clock_I (.I(clknet_5_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_121_clock_I (.I(clknet_5_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_120_clock_I (.I(clknet_5_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_119_clock_I (.I(clknet_5_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_118_clock_I (.I(clknet_5_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_309_clock_I (.I(clknet_5_16_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13393__CLK (.I(clknet_5_16_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_307_clock_I (.I(clknet_5_16_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_306_clock_I (.I(clknet_5_16_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_305_clock_I (.I(clknet_5_16_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_304_clock_I (.I(clknet_5_16_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_303_clock_I (.I(clknet_5_16_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_302_clock_I (.I(clknet_5_16_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_301_clock_I (.I(clknet_5_16_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_312_clock_I (.I(clknet_5_17_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_311_clock_I (.I(clknet_5_17_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_310_clock_I (.I(clknet_5_17_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_300_clock_I (.I(clknet_5_17_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_299_clock_I (.I(clknet_5_17_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_298_clock_I (.I(clknet_5_17_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_297_clock_I (.I(clknet_5_17_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_296_clock_I (.I(clknet_5_17_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_295_clock_I (.I(clknet_5_17_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_323_clock_I (.I(clknet_5_18_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_322_clock_I (.I(clknet_5_18_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_321_clock_I (.I(clknet_5_18_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_320_clock_I (.I(clknet_5_18_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_319_clock_I (.I(clknet_5_18_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_318_clock_I (.I(clknet_5_18_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_317_clock_I (.I(clknet_5_18_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_316_clock_I (.I(clknet_5_18_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_315_clock_I (.I(clknet_5_18_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_235_clock_I (.I(clknet_5_18_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_234_clock_I (.I(clknet_5_18_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_233_clock_I (.I(clknet_5_18_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_314_clock_I (.I(clknet_5_19_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_313_clock_I (.I(clknet_5_19_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_244_clock_I (.I(clknet_5_19_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_243_clock_I (.I(clknet_5_19_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_242_clock_I (.I(clknet_5_19_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_241_clock_I (.I(clknet_5_19_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_240_clock_I (.I(clknet_5_19_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_239_clock_I (.I(clknet_5_19_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_238_clock_I (.I(clknet_5_19_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_237_clock_I (.I(clknet_5_19_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_236_clock_I (.I(clknet_5_19_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_294_clock_I (.I(clknet_5_20_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_293_clock_I (.I(clknet_5_20_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_292_clock_I (.I(clknet_5_20_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_291_clock_I (.I(clknet_5_20_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_290_clock_I (.I(clknet_5_20_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_289_clock_I (.I(clknet_5_20_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_288_clock_I (.I(clknet_5_20_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_287_clock_I (.I(clknet_5_20_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_286_clock_I (.I(clknet_5_20_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_285_clock_I (.I(clknet_5_20_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_272_clock_I (.I(clknet_5_20_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_271_clock_I (.I(clknet_5_20_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_270_clock_I (.I(clknet_5_20_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_284_clock_I (.I(clknet_5_21_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_283_clock_I (.I(clknet_5_21_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_282_clock_I (.I(clknet_5_21_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_281_clock_I (.I(clknet_5_21_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_280_clock_I (.I(clknet_5_21_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_279_clock_I (.I(clknet_5_21_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_278_clock_I (.I(clknet_5_21_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_277_clock_I (.I(clknet_5_21_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_276_clock_I (.I(clknet_5_21_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_275_clock_I (.I(clknet_5_21_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_274_clock_I (.I(clknet_5_21_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_273_clock_I (.I(clknet_5_21_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_269_clock_I (.I(clknet_5_22_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_268_clock_I (.I(clknet_5_22_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_267_clock_I (.I(clknet_5_22_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_253_clock_I (.I(clknet_5_22_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_252_clock_I (.I(clknet_5_22_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_251_clock_I (.I(clknet_5_22_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_250_clock_I (.I(clknet_5_22_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_249_clock_I (.I(clknet_5_22_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_248_clock_I (.I(clknet_5_22_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13115__CLK (.I(clknet_5_22_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_246_clock_I (.I(clknet_5_22_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_245_clock_I (.I(clknet_5_22_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_266_clock_I (.I(clknet_5_23_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_265_clock_I (.I(clknet_5_23_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_264_clock_I (.I(clknet_5_23_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_263_clock_I (.I(clknet_5_23_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_262_clock_I (.I(clknet_5_23_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_261_clock_I (.I(clknet_5_23_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_260_clock_I (.I(clknet_5_23_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_259_clock_I (.I(clknet_5_23_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_258_clock_I (.I(clknet_5_23_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_257_clock_I (.I(clknet_5_23_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_256_clock_I (.I(clknet_5_23_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_255_clock_I (.I(clknet_5_23_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_254_clock_I (.I(clknet_5_23_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_232_clock_I (.I(clknet_5_24_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_231_clock_I (.I(clknet_5_24_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_230_clock_I (.I(clknet_5_24_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_149_clock_I (.I(clknet_5_24_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_148_clock_I (.I(clknet_5_24_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_147_clock_I (.I(clknet_5_24_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_146_clock_I (.I(clknet_5_24_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_145_clock_I (.I(clknet_5_24_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_144_clock_I (.I(clknet_5_24_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_143_clock_I (.I(clknet_5_24_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_229_clock_I (.I(clknet_5_25_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_228_clock_I (.I(clknet_5_25_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_227_clock_I (.I(clknet_5_25_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_226_clock_I (.I(clknet_5_25_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_225_clock_I (.I(clknet_5_25_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_224_clock_I (.I(clknet_5_25_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_223_clock_I (.I(clknet_5_25_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_153_clock_I (.I(clknet_5_25_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_152_clock_I (.I(clknet_5_25_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_151_clock_I (.I(clknet_5_25_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_150_clock_I (.I(clknet_5_25_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_167_clock_I (.I(clknet_5_26_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_166_clock_I (.I(clknet_5_26_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_165_clock_I (.I(clknet_5_26_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_164_clock_I (.I(clknet_5_26_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_163_clock_I (.I(clknet_5_26_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_162_clock_I (.I(clknet_5_26_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_161_clock_I (.I(clknet_5_26_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_160_clock_I (.I(clknet_5_26_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_159_clock_I (.I(clknet_5_26_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_158_clock_I (.I(clknet_5_26_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_157_clock_I (.I(clknet_5_26_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_156_clock_I (.I(clknet_5_26_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_184_clock_I (.I(clknet_5_27_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_182_clock_I (.I(clknet_5_27_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_177_clock_I (.I(clknet_5_27_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12690__CLK (.I(clknet_5_27_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_175_clock_I (.I(clknet_5_27_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_174_clock_I (.I(clknet_5_27_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_173_clock_I (.I(clknet_5_27_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_172_clock_I (.I(clknet_5_27_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_171_clock_I (.I(clknet_5_27_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_170_clock_I (.I(clknet_5_27_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_169_clock_I (.I(clknet_5_27_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_168_clock_I (.I(clknet_5_27_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_155_clock_I (.I(clknet_5_27_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_154_clock_I (.I(clknet_5_27_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_222_clock_I (.I(clknet_5_28_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_221_clock_I (.I(clknet_5_28_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_220_clock_I (.I(clknet_5_28_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_219_clock_I (.I(clknet_5_28_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_218_clock_I (.I(clknet_5_28_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_217_clock_I (.I(clknet_5_28_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_216_clock_I (.I(clknet_5_28_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_215_clock_I (.I(clknet_5_28_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_214_clock_I (.I(clknet_5_28_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_201_clock_I (.I(clknet_5_28_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_200_clock_I (.I(clknet_5_28_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_199_clock_I (.I(clknet_5_28_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_213_clock_I (.I(clknet_5_29_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_212_clock_I (.I(clknet_5_29_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_211_clock_I (.I(clknet_5_29_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_210_clock_I (.I(clknet_5_29_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_209_clock_I (.I(clknet_5_29_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_208_clock_I (.I(clknet_5_29_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_207_clock_I (.I(clknet_5_29_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_206_clock_I (.I(clknet_5_29_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_205_clock_I (.I(clknet_5_29_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_204_clock_I (.I(clknet_5_29_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_203_clock_I (.I(clknet_5_29_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_202_clock_I (.I(clknet_5_29_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_198_clock_I (.I(clknet_5_30_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_197_clock_I (.I(clknet_5_30_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_185_clock_I (.I(clknet_5_30_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_183_clock_I (.I(clknet_5_30_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_181_clock_I (.I(clknet_5_30_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_180_clock_I (.I(clknet_5_30_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_179_clock_I (.I(clknet_5_30_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_178_clock_I (.I(clknet_5_30_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_196_clock_I (.I(clknet_5_31_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_195_clock_I (.I(clknet_5_31_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_194_clock_I (.I(clknet_5_31_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_193_clock_I (.I(clknet_5_31_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_192_clock_I (.I(clknet_5_31_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_191_clock_I (.I(clknet_5_31_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_190_clock_I (.I(clknet_5_31_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_189_clock_I (.I(clknet_5_31_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_188_clock_I (.I(clknet_5_31_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_187_clock_I (.I(clknet_5_31_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_186_clock_I (.I(clknet_5_31_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_3__f_clock_a_I (.I(clknet_0_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_2__f_clock_a_I (.I(clknet_0_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_1__f_clock_a_I (.I(clknet_0_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_0__f_clock_a_I (.I(clknet_0_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12009__CLK (.I(clknet_2_0__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12013__CLK (.I(clknet_2_0__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12027__CLK (.I(clknet_2_0__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12037__CLK (.I(clknet_2_0__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12051__CLK (.I(clknet_2_0__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12053__CLK (.I(clknet_2_0__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12061__CLK (.I(clknet_2_0__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12069__CLK (.I(clknet_2_0__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12089__CLK (.I(clknet_2_0__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12011__CLK (.I(clknet_2_1__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12021__CLK (.I(clknet_2_1__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12023__CLK (.I(clknet_2_1__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12057__CLK (.I(clknet_2_1__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12059__CLK (.I(clknet_2_1__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12067__CLK (.I(clknet_2_1__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12071__CLK (.I(clknet_2_1__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12073__CLK (.I(clknet_2_1__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12079__CLK (.I(clknet_2_1__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12087__CLK (.I(clknet_2_1__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12007__CLK (.I(clknet_2_2__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12015__CLK (.I(clknet_2_2__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12017__CLK (.I(clknet_2_2__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12019__CLK (.I(clknet_2_2__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12029__CLK (.I(clknet_2_2__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12039__CLK (.I(clknet_2_2__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12043__CLK (.I(clknet_2_2__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12045__CLK (.I(clknet_2_2__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12047__CLK (.I(clknet_2_2__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12055__CLK (.I(clknet_2_2__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12075__CLK (.I(clknet_2_2__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12077__CLK (.I(clknet_2_2__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12085__CLK (.I(clknet_2_2__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12005__CLK (.I(clknet_2_3__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12025__CLK (.I(clknet_2_3__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12031__CLK (.I(clknet_2_3__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12033__CLK (.I(clknet_2_3__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12035__CLK (.I(clknet_2_3__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12041__CLK (.I(clknet_2_3__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12049__CLK (.I(clknet_2_3__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12063__CLK (.I(clknet_2_3__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12065__CLK (.I(clknet_2_3__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12091__CLK (.I(clknet_2_3__leaf_clock_a));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12081__D (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1577 ();
endmodule

