* NGSPICE file created from user_proj_example.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

.subckt user_proj_example io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ irq[0] irq[1] irq[2] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102]
+ la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107]
+ la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112]
+ la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117]
+ la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122]
+ la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127]
+ la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17]
+ la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22]
+ la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28]
+ la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33]
+ la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39]
+ la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44]
+ la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4]
+ la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60]
+ la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66]
+ la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71]
+ la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77]
+ la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82]
+ la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88]
+ la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93]
+ la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99]
+ la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XFILLER_95_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input108_I wbs_we_i vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input73_I wbs_dat_i[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__429__I _123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_501_ _199_ _202_ _014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_432_ _133_ _134_ net93 _138_ _145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_2589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__760__CLK clknet_3_6__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_363_ net35 _071_ _078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__568__A1 net162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__559__A1 _247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__495__C2 net74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_415_ net146 _130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput231 net231 wbs_dat_o[28] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput242 net242 wbs_dat_o[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput220 net220 wbs_dat_o[18] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_138_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input36_I la_oenb[33] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__442__I net172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_895_ net138 net129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__352__I net210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_680_ _338_ _057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__900__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_878_ net138 net111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__392__A2 _106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__604__C2 net92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__604__B1 _256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__383__A2 _091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__717__CLK clknet_3_4__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_732_ _036_ clknet_3_1__leaf_counter.clk net236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_663_ net219 net154 _321_ _329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_594_ net28 _282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__374__A2 _078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_715_ _019_ clknet_3_7__leaf_counter.clk net155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_76_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_646_ net212 _304_ _319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_577_ _256_ _267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__595__A2 _282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__360__I _075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input66_I la_oenb[63] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_500_ net14 _099_ _175_ _201_ _194_ net75 _202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA_output222_I net222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_431_ _142_ _127_ _143_ _144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_362_ _065_ _077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_629_ net233 net168 _309_ _310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output172_I net172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__495__A1 net13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_414_ _128_ _129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__903__I net146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_7__f_counter.clk clknet_0_counter.clk clknet_3_7__leaf_counter.clk vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput210 net210 wbs_ack_o vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput221 net221 wbs_dat_o[19] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput232 net232 wbs_dat_o[29] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__477__A1 net177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__750__CLK clknet_3_2__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input29_I la_data_in[60] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__401__A1 _112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__468__A1 _123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_894_ net138 net128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__402__B _106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_877_ net138 net110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__628__I _308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__604__A1 net30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input96_I wbs_dat_i[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__383__A3 _092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_731_ _035_ clknet_3_0__leaf_counter.clk net233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_662_ _328_ _049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_593_ _267_ _280_ _281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__374__A3 _088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__911__I net176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_929_ net164 net196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input11_I la_data_in[42] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_714_ _018_ clknet_3_4__leaf_counter.clk net154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_645_ _318_ _042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_576_ net161 net162 _251_ _266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__595__A3 _072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__906__I net171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input3_I la_data_in[34] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__707__CLK clknet_3_6__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input59_I la_oenb[56] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output215_I net215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_430_ _136_ _130_ net168 _143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_361_ _076_ _000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_628_ _308_ _309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_127_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_559_ _247_ _243_ _251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__371__I _085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output165_I net165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__495__A2 _102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_413_ _123_ _127_ _128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput200 net200 la_data_out[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_47_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput222 net222 wbs_dat_o[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput233 net233 wbs_dat_o[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput211 net211 wbs_dat_o[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__477__A2 net176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__401__A2 _113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_893_ net138 net127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__640__A2 _304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__914__I net148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input41_I la_oenb[38] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__622__A2 _304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_876_ net138 net145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__909__I net174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__377__A1 net46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__740__CLK clknet_3_0__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__554__I net160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__383__A4 _097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input89_I wbs_dat_i[26] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__540__A1 _231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_730_ _034_ clknet_3_1__leaf_counter.clk net222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_661_ net218 net153 _321_ _328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_592_ _275_ _271_ _278_ _280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_928_ net163 net195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__598__A1 net63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__696__D _000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__589__A1 _274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput100 wbs_dat_i[7] net100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_713_ _017_ clknet_3_4__leaf_counter.clk net153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__459__I net175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_644_ net242 net177 _314_ _318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_575_ net163 _265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__922__I net156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__504__A1 _203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_360_ _075_ _076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__917__I net151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_627_ _074_ _308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_558_ net58 _165_ _250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_489_ net148 _192_ _193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_9_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input106_I wbs_sel_i[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input71_I wbs_dat_i[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output158_I net158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_412_ _124_ _126_ _127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput201 net201 la_data_out[30] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_12_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput234 net234 wbs_dat_o[30] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput212 net212 wbs_dat_o[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput223 net223 wbs_dat_o[20] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_114_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__401__A3 _114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_892_ net138 net126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__930__I net165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__395__A2 _109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_3__f_counter.clk clknet_0_counter.clk clknet_3_3__leaf_counter.clk vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_115_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input34_I la_data_in[65] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_875_ net138 net144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__925__I net160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__688__I0 net231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__368__A2 _082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__570__I _260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__679__I0 net227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_660_ _210_ _324_ _327_ _048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_591_ net164 _278_ _270_ _279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_16_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_927_ net162 net194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__655__I _076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__513__A2 _212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput101 wbs_dat_i[8] net101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__730__CLK clknet_3_1__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_712_ _016_ clknet_3_7__leaf_counter.clk net152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_643_ _317_ _041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_574_ _260_ _264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__753__CLK clknet_3_6__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__498__A1 net149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_626_ _307_ _034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_557_ _246_ _249_ _023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_488_ _191_ _167_ _169_ _183_ _192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__933__I net169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__489__A1 net148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__413__A1 _123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input64_I la_oenb[61] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output220_I net220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_411_ _125_ net103 _126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__928__I net163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_609_ net169 _294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput235 net235 wbs_dat_o[31] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput213 net213 wbs_dat_o[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput224 net224 wbs_dat_o[21] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput202 net202 la_data_out[31] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_126_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__401__A4 _115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output170_I net170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_891_ net138 net125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__684__S _337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__561__B1 _216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__561__C2 net86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__616__A1 _292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__658__I _075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input27_I la_data_in[58] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__679__S _337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_874_ net138 net143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__688__I1 net166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__679__I1 net162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_590_ net165 _278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_926_ net161 net193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__620__B _188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input94_I wbs_dat_i[30] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput102 wbs_dat_i[9] net102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_711_ _015_ clknet_3_7__leaf_counter.clk net151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_642_ net241 net176 _314_ _317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_573_ net60 _151_ _263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_909_ net174 net206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__431__A2 _127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_625_ net222 _136_ _306_ _307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_556_ net23 _107_ _216_ _248_ _233_ net85 _249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_17_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_487_ net147 _191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_13_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I la_data_in[32] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__413__A2 _127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__720__CLK clknet_3_7__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input57_I la_oenb[54] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__404__A2 net66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_410_ net108 _125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_608_ _275_ _278_ net166 _271_ _293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_17_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__743__CLK clknet_3_1__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_539_ _231_ net156 _228_ _235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_18_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput214 net214 wbs_dat_o[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput225 net225 wbs_dat_o[22] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput203 net203 la_data_out[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput236 net236 wbs_dat_o[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_142_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output163_I net163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_890_ net138 net124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__389__A1 _099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__561__A1 net24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__616__A2 _294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_873_ net138 net142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__516__A1 _138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_925_ net160 net192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input87_I wbs_dat_i[24] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput103 wbs_sel_i[0] net103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_710_ _014_ clknet_3_7__leaf_counter.clk net150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_131_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_641_ _168_ _000_ _316_ _040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_572_ _246_ _262_ _025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_908_ net173 net205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_0 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_624_ _074_ _306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_555_ _247_ _243_ _248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_486_ _172_ _190_ _011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__497__I _077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__651__I0 net214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_607_ net167 _292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_538_ _223_ _234_ _019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_469_ _175_ _176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput215 net215 wbs_dat_o[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput226 net226 wbs_dat_o[23] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput204 net204 la_data_out[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_114_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput237 net237 wbs_dat_o[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_4_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__398__A2 _106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__642__I0 net241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input104_I wbs_sel_i[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__870__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output156_I net156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__389__A2 _100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__561__A2 _250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__710__CLK clknet_3_7__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__733__CLK clknet_3_1__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_872_ net138 net141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__470__A1 _168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__756__CLK clknet_3_6__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input32_I la_data_in[63] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__461__A1 net174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__516__A2 _214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_924_ net159 net191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_340 la_data_out[119] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_144_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__691__A1 _292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__443__A1 net171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput104 wbs_sel_i[1] net104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_640_ net240 _304_ _316_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__434__A1 net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_571_ net25 _081_ _257_ _259_ _261_ net87 _262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_17_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_2__f_counter.clk_I clknet_0_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_907_ net172 net204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__873__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_623_ _131_ _000_ _305_ _033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_554_ net160 _247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_60_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_485_ net11 _100_ _176_ _189_ _180_ net72 _190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_129_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__868__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__552__B _188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_606_ net167 net169 _288_ _291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_537_ net19 _114_ _217_ _232_ _233_ net80 _234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__651__I1 net149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_468_ _123_ _174_ _175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_399_ net53 _109_ _114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput205 net205 la_data_out[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput216 net216 wbs_dat_o[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_12_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput238 net238 wbs_dat_o[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput227 net227 wbs_dat_o[24] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_5_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__619__A1 net32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__619__B2 net95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__642__I1 net176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input62_I la_oenb[59] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output149_I net149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__389__A3 _102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__633__I1 _153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_7__f_counter.clk_I clknet_0_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__537__C2 net80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__881__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_871_ net138 net140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__470__A2 _169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__876__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input25_I la_data_in[56] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__461__A2 net173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__700__CLK clknet_3_3__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_923_ net158 net190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_330 la_data_out[109] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_341 la_data_out[120] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__691__A2 _339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__443__A2 net168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__723__CLK clknet_3_5__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput105 wbs_sel_i[2] net105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__682__A2 _326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_570_ _260_ _261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_906_ net171 net203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__746__CLK clknet_3_2__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_699_ _003_ clknet_3_3__leaf_counter.clk net168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input92_I wbs_dat_i[29] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_622_ net211 _304_ _305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_553_ _066_ _246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_484_ net147 _184_ _189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_13_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__591__A1 net164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__646__A2 _304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__582__A1 _265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__884__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__573__A1 net60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_605_ _274_ _290_ _030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_536_ _220_ _233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_467_ _124_ _173_ _174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__564__A1 _124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_398_ net38 _106_ _113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput217 net217 wbs_dat_o[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput206 net206 la_data_out[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_126_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput239 net239 wbs_dat_o[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput228 net228 wbs_dat_o[25] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_5_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__619__A2 _302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__555__A1 _247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__879__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input55_I la_oenb[52] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__491__C2 net73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__389__A4 _103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_519_ _210_ _205_ _218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__537__A1 net19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__528__A1 net153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output161_I net161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_870_ net138 net139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__519__A1 _210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__455__B1 _128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__455__C2 net99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__461__A3 net172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input18_I la_data_in[49] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__892__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_922_ net156 net188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__437__B1 _129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_320 la_data_out[99] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_11_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_342 la_data_out[121] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_331 la_data_out[110] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__443__A3 net157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__600__B1 _256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__600__C2 net91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__887__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput106 wbs_sel_i[3] net106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__698__CLK clknet_3_2__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_905_ net168 net200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__425__A3 net82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_698_ _002_ clknet_3_2__leaf_counter.clk net157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__672__I0 net224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input85_I wbs_dat_i[22] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output241_I net241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__410__I net108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_621_ _075_ _304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__663__I0 net219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_552_ _244_ _245_ _188_ _022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_483_ _186_ _187_ _188_ _010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_13_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__591__A2 _278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__713__CLK clknet_3_4__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__476__B net177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__736__CLK clknet_3_0__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_604_ net30 _093_ _256_ _289_ _261_ net92 _290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_2863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_535_ _231_ _228_ _232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_33_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_466_ net108 net104 _173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_397_ net52 _101_ _112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__564__A2 _254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput207 net207 la_data_out[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_138_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput218 net218 wbs_dat_o[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput229 net229 wbs_dat_o[26] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_4_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__759__CLK clknet_3_3__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input48_I la_oenb[45] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__895__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__491__A1 net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_518_ _216_ _217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_449_ _153_ _154_ _159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__537__A2 _114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input102_I wbs_dat_i[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__528__A2 net154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output154_I net154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__455__A1 net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_921_ net155 net187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__437__A1 net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_321 la_data_out[100] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_310 la_data_out[89] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_proj_example_343 la_data_out[122] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_332 la_data_out[111] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__428__A1 net168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__443__A4 net146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__600__A1 net29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput107 wbs_stb_i net107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input30_I la_data_in[61] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_904_ net157 net189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__425__A4 _138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_697_ _001_ clknet_3_0__leaf_counter.clk net146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__672__I1 net159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input78_I wbs_dat_i[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__898__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_620_ _301_ _303_ _188_ _032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__407__A4 _121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_551_ net22 _105_ _221_ net84 _245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__663__I1 net154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_482_ _065_ _188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__500__C2 net75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_749_ _053_ clknet_3_2__leaf_counter.clk net223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_603_ net167 _288_ _289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_534_ net155 _231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_465_ _077_ _172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_396_ _105_ _107_ _108_ _110_ _111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_13_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput208 net208 la_data_out[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_114_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput219 net219 wbs_dat_o[17] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_141_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__491__A2 _092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__416__I _130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__703__CLK clknet_3_3__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_517_ _142_ _215_ _216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_448_ _150_ _158_ _005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_379_ net61 _079_ _094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__726__CLK clknet_3_5__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input60_I la_oenb[57] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output147_I net147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__347__S net68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__455__A2 _115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__749__CLK clknet_3_2__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__694__A2 _306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__446__A2 _126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_920_ net154 net186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__437__A2 _113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_311 la_data_out[90] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_300 la_data_out[79] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xuser_proj_example_344 la_data_out[123] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_333 la_data_out[112] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_322 la_data_out[101] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__676__A2 _326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__428__A2 _136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_6__f_counter.clk clknet_0_counter.clk clknet_3_6__leaf_counter.clk vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_53_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput108 wbs_we_i net108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input23_I la_data_in[54] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__625__S _306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__424__I _124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_903_ net146 net178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_696_ _000_ clknet_3_1__leaf_counter.clk net210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput90 wbs_dat_i[27] net90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output227_I net227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_550_ net159 _241_ _243_ _217_ _244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_17_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__419__I net103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_481_ net10 _103_ _180_ net102 _187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__576__A1 net161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__500__A1 net14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_748_ _052_ clknet_3_2__leaf_counter.clk net221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_679_ net227 net162 _337_ _338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__567__A1 net161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__558__A1 net58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input90_I wbs_dat_i[27] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output177_I net177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_602_ net164 net165 net166 _270_ _288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_2821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_533_ _223_ _230_ _018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_464_ _150_ _171_ _008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__549__A1 net155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_395_ net40 _109_ _110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput209 net209 la_data_out[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_5_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__485__C2 net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__522__I _220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_516_ _138_ _214_ _215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__607__I net167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_447_ net5 _152_ _129_ _155_ _157_ net97 _158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_378_ net64 _079_ _093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input53_I la_oenb[50] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_312 la_data_out[91] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_301 la_data_out[80] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__373__A2 _071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_345 la_data_out[124] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_334 la_data_out[113] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_323 la_data_out[102] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__716__CLK clknet_3_4__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__428__A3 _130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input16_I la_data_in[47] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__739__CLK clknet_3_0__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__440__I _072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_902_ net138 net137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__666__I0 net220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_695_ _299_ _339_ _346_ _064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__615__I net170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input8_I la_data_in[39] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__525__I _066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput91 wbs_dat_i[28] net91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput80 wbs_dat_i[18] net80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_480_ _176_ _185_ _186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__576__A2 net162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__500__A2 _099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_747_ _051_ clknet_3_2__leaf_counter.clk net220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_678_ _075_ _337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_95_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input83_I wbs_dat_i[20] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__494__A1 net149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_601_ _274_ _287_ _029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_532_ net18 _112_ _221_ net79 _229_ _230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_144_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_463_ net8 _166_ _128_ _170_ _157_ net100 _171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__549__A2 net156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_394_ _085_ _109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__485__A1 net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__476__A1 net176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__467__A1 _124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_515_ net105 _125_ _214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_446_ _156_ _126_ _157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_377_ net46 _080_ _092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__449__A1 _153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input46_I la_oenb[43] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__612__B2 net94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__612__A1 net31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_429_ _123_ _142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput1 la_data_in[32] net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__603__A1 net167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input100_I wbs_dat_i[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output152_I net152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_302 la_data_out[81] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_11_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_346 la_data_out[125] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_335 la_data_out[114] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_324 la_data_out[103] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_313 la_data_out[92] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__901__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__684__I1 _275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__348__I _065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__588__C2 net89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__512__C2 net77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_901_ net138 net136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput190 net190 la_data_out[20] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_134_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__666__I1 _231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__596__C _283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_694_ net235 _306_ _346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput81 wbs_dat_i[19] net81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput70 wbs_cyc_i net70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_3_2__f_counter.clk clknet_0_counter.clk clknet_3_2__leaf_counter.clk vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_118_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput92 wbs_dat_i[29] net92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__648__I1 net148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__706__CLK clknet_3_7__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_746_ _050_ clknet_3_2__leaf_counter.clk net219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_677_ _268_ _324_ _336_ _056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__361__I _076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__729__CLK clknet_3_1__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__536__I _220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input76_I wbs_dat_i[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output232_I net232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_600_ net29 _285_ _256_ _286_ _261_ net91 _287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_3524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_531_ _224_ _225_ _228_ _229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_2_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_462_ _168_ _169_ _170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_393_ net55 _106_ _108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__485__A2 _100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_729_ _033_ clknet_3_1__leaf_counter.clk net211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__356__I _071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__467__A2 _173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_514_ net51 _165_ _213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_445_ _073_ _156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_376_ net54 _086_ _091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__904__I net157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input39_I la_oenb[36] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__385__A1 net45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_428_ net168 _136_ _130_ _141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__376__A1 net54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_359_ _074_ _075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput2 la_data_in[33] net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__603__A2 _288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__358__A1 _065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_303 la_data_out[82] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_336 la_data_out[115] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_325 la_data_out[104] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_314 la_data_out[93] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_137_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_347 la_data_out[126] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_13_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__597__A1 _274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__364__I _069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__588__A1 net27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__512__A1 net16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_900_ net138 net135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput191 net191 la_data_out[21] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput180 net180 la_data_out[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_87_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_0__f_counter.clk_I clknet_0_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_693_ _294_ _339_ _345_ _063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__579__A1 net162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__912__I net177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__503__A1 net150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__359__I _074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput82 wbs_dat_i[1] net82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput71 wbs_dat_i[0] net71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput60 la_oenb[57] net60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput93 wbs_dat_i[2] net93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input21_I la_data_in[52] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_745_ _049_ clknet_3_0__leaf_counter.clk net218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_676_ net226 _326_ _336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__907__I net172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input69_I wb_rst_i vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_530_ _227_ _228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output225_I net225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_461_ net174 net173 net172 _154_ _169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_57_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_392_ net57 _106_ _107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__637__I _308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_728_ _032_ clknet_3_7__leaf_counter.clk net170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_659_ net217 _326_ _327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output175_I net175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_5__f_counter.clk_I clknet_0_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__457__I _072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_513_ _199_ _212_ _016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_444_ _153_ _154_ _155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_375_ net43 _080_ _090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__719__CLK clknet_3_7__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__920__I net154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__915__I net149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_427_ net138 _140_ _002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_358_ _065_ _073_ _074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__650__I _308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput3 la_data_in[34] net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input51_I la_oenb[48] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output138_I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_337 la_data_out[116] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_326 la_data_out[105] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_315 la_data_out[94] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_304 la_data_out[83] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_11_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_348 la_data_out[127] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__521__A2 _214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input99_I wbs_dat_i[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__512__A2 _118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput170 net170 io_out[31] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_133_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput181 net181 la_data_out[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput192 net192 la_data_out[22] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_692_ net234 _306_ _345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__579__A2 net163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__465__I _077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__503__A2 net149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput72 wbs_dat_i[10] net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput50 la_oenb[47] net50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput61 la_oenb[58] net61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput83 wbs_dat_i[20] net83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput94 wbs_dat_i[30] net94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input14_I la_data_in[45] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__430__A1 _136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__752__CLK clknet_3_1__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_744_ _048_ clknet_3_0__leaf_counter.clk net217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_675_ _247_ _324_ _335_ _055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__421__A1 _077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__923__I net158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__488__A1 _191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I la_data_in[37] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__660__A1 _210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__412__A1 _124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_460_ _167_ _168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_391_ _085_ _106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__918__I net152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_727_ _031_ clknet_3_7__leaf_counter.clk net169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_658_ _075_ _326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_589_ _274_ _277_ _027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input81_I wbs_dat_i[19] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output168_I net168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_512_ net16 _118_ _175_ _211_ _194_ net77 _212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_2688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_443_ net171 net168 net157 net146 _154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_2_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_374_ _087_ _078_ _088_ _089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_13_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__551__B1 _221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__606__A1 net167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__542__B1 _221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_426_ net2 _088_ _129_ _137_ _139_ _140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_14_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_357_ _068_ _072_ _073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__931__I net166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 la_data_in[35] net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input44_I la_oenb[41] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__709__CLK clknet_3_6__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_327 la_data_out[106] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_316 la_data_out[95] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_305 la_data_out[84] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_11_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_338 la_data_out[117] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_139_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__926__I net161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_409_ _087_ _124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__610__B _294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput160 net160 io_out[22] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output150_I net150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput171 net171 io_out[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_82_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput182 net182 la_data_out[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput193 net193 la_data_out[23] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_88_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_760_ _064_ clknet_3_6__leaf_counter.clk net235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_691_ _292_ _339_ _344_ _062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__503__A3 net148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__430__B net168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_889_ net138 net123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__391__I _085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput40 la_oenb[37] net40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput51 la_oenb[48] net51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput62 la_oenb[59] net62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput73 wbs_dat_i[11] net73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput95 wbs_dat_i[31] net95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput84 wbs_dat_i[21] net84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__566__I _256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__430__A2 _130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_743_ _047_ clknet_3_1__leaf_counter.clk net216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_674_ net225 _326_ _335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__660__A2 _324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__386__I _085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__412__A2 _126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__403__A2 _109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_390_ net56 _101_ _105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_726_ _030_ clknet_3_5__leaf_counter.clk net167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_91_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_657_ _203_ _324_ _325_ _047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_588_ net27 _094_ _257_ _276_ _261_ net89 _277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_16_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__934__I net170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__742__CLK clknet_3_2__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input74_I wbs_dat_i[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output230_I net230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_511_ _210_ _205_ _211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_442_ net172 _153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_373_ net36 _071_ _088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__560__A1 net161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__929__I net164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_709_ _013_ clknet_3_6__leaf_counter.clk net149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__379__A1 net61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__613__B _188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__551__B2 net84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__551__A1 net22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__606__A2 net169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__574__I _260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__542__B2 net81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__542__A1 net20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_425_ _133_ _134_ net82 _138_ _139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_14_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_356_ _071_ _072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput5 la_data_in[36] net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__394__I _085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input37_I la_oenb[34] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_328 la_data_out[107] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_317 la_data_out[96] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_306 la_data_out[85] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__515__A1 net105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_339 la_data_out[118] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_13_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__451__C2 net98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__451__B1 _128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_408_ _084_ _089_ _098_ _122_ _123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_119_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput161 net161 io_out[23] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput150 net150 io_out[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput172 net172 io_out[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_121_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput183 net183 la_data_out[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput194 net194 la_data_out[24] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_101_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_690_ net232 _306_ _344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__433__B1 _141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_888_ net138 net122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput30 la_data_in[61] net30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput63 la_oenb[60] net63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput41 la_oenb[38] net41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput52 la_oenb[49] net52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput74 wbs_dat_i[12] net74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput96 wbs_dat_i[3] net96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput85 wbs_dat_i[22] net85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_742_ _046_ clknet_3_2__leaf_counter.clk net215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_673_ _334_ _054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__488__A3 _169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__616__B _299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__577__I _256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__688__S _337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__487__I net147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_725_ _029_ clknet_3_4__leaf_counter.clk net166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_90_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_656_ net216 _304_ _325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_587_ _275_ _271_ _276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_16_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__397__A2 _101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input67_I la_oenb[64] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_510_ net152 _210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_3369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_441_ net39 _151_ _152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__388__A2 _101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_372_ _068_ _086_ _087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_13_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_708_ _012_ clknet_3_6__leaf_counter.clk net148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_17_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_639_ _315_ _039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__551__A2 _105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__606__A3 _288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__590__I net165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__542__A2 _091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output173_I net173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_424_ _124_ _138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_355_ _070_ _071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__433__C _145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__732__CLK clknet_3_1__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput6 la_data_in[37] net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__585__I _066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_318 la_data_out[97] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_307 la_data_out[86] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__515__A2 _125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_329 la_data_out[108] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_137_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__755__CLK clknet_3_2__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__451__A1 net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_407_ _104_ _111_ _116_ _121_ _122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_30_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__690__A1 net232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput151 net151 io_out[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput140 net140 io_oeb[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_88_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput173 net173 io_out[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput162 net162 io_out[24] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_115_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput184 net184 la_data_out[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput195 net195 la_data_out[25] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__433__A1 net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_887_ net138 net121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput31 la_data_in[62] net31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput20 la_data_in[51] net20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput64 la_oenb[61] net64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput42 la_oenb[39] net42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput53 la_oenb[50] net53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput86 wbs_dat_i[23] net86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput97 wbs_dat_i[4] net97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput75 wbs_dat_i[13] net75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input97_I wbs_dat_i[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_741_ _045_ clknet_3_2__leaf_counter.clk net214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_672_ net224 net159 _330_ _334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input12_I la_data_in[43] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_724_ _028_ clknet_3_5__leaf_counter.clk net165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_655_ _076_ _324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_586_ net164 _275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__618__A1 net66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__678__I _075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input4_I la_data_in[35] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_440_ _072_ _151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_371_ _085_ _086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__545__C2 net83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_707_ _011_ clknet_3_6__leaf_counter.clk net147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_638_ net239 net174 _314_ _315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_569_ _156_ _254_ _260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__871__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output166_I net166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_423_ _136_ _130_ _137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_354_ _069_ _070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput7 la_data_in[38] net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xuser_proj_example_319 la_data_out[98] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_308 la_data_out[87] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_136_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__451__A2 _110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_406_ _117_ _118_ _119_ _120_ _121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_109_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__690__A2 _306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput130 net130 io_oeb[29] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput152 net152 io_out[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput141 net141 io_oeb[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_86_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput163 net163 io_out[25] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput174 net174 io_out[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_134_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput185 net185 la_data_out[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA_input42_I la_oenb[39] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput196 net196 la_data_out[26] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_88_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__433__A2 _082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__722__CLK clknet_3_5__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_886_ net138 net119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput10 la_data_in[41] net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 la_data_in[52] net21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput32 la_data_in[63] net32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput43 la_oenb[40] net43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput54 la_oenb[51] net54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput98 wbs_dat_i[5] net98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput76 wbs_dat_i[14] net76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput65 la_oenb[62] net65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput87 wbs_dat_i[24] net87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__745__CLK clknet_3_0__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_740_ _044_ clknet_3_0__leaf_counter.clk net213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__406__A2 _118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_671_ _333_ _053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_869_ net138 net131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__874__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__572__A1 _246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_723_ _027_ clknet_3_5__leaf_counter.clk net164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_654_ _323_ _046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_585_ _066_ _274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__563__A1 _125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__869__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_370_ _069_ _085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__545__A1 net21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_706_ _010_ clknet_3_7__leaf_counter.clk net177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_637_ _308_ _314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_568_ net162 _258_ _259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_17_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_499_ net150 _200_ _201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_125_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input107_I wbs_stb_i vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__527__A1 net153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input72_I wbs_dat_i[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output159_I net159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__463__C2 net100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__463__B1 _128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_422_ net157 _136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_353_ net107 net70 _069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_126_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput8 la_data_in[39] net8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__882__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_309 la_data_out[88] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_11_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_405_ net42 net51 _070_ _120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput142 net142 io_oeb[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput120 net120 io_oeb[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput131 net131 io_oeb[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput164 net164 io_out[26] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput153 net153 io_out[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput175 net175 io_out[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_82_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput186 net186 la_data_out[17] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__877__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput197 net197 la_data_out[27] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_101_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input35_I la_oenb[32] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_885_ net138 net118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput11 la_data_in[42] net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 la_data_in[53] net22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__697__CLK clknet_3_0__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput33 la_data_in[64] net33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput44 la_oenb[41] net44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput55 la_oenb[52] net55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput77 wbs_dat_i[15] net77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput66 la_oenb[63] net66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput88 wbs_dat_i[25] net88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput99 wbs_dat_i[6] net99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output239_I net239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_670_ net223 net158 _330_ _333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_868_ net138 net120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__653__I0 net215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__712__CLK clknet_3_7__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__890__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_722_ _026_ clknet_3_5__leaf_counter.clk net163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_653_ net215 net150 _321_ _323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_584_ _246_ _273_ _026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__735__CLK clknet_3_2__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_5__f_counter.clk clknet_0_counter.clk clknet_3_5__leaf_counter.clk vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__885__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__545__A2 _108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__758__CLK clknet_3_3__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__481__A1 net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_705_ _009_ clknet_3_6__leaf_counter.clk net176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__481__B2 net102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_636_ _313_ _038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_567_ net161 _251_ _258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_498_ net149 _196_ _200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input65_I la_oenb[62] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__463__A1 net8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output221_I net221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_421_ _077_ _132_ _135_ _001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_352_ net210 _068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__454__A1 net174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 la_data_in[40] net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_619_ net32 _302_ _264_ net95 _303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__693__A1 _294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output171_I net171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_404_ net49 net66 _109_ _119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_127_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__675__A1 _247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__427__A1 net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput110 net110 io_oeb[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_133_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput132 net132 io_oeb[30] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput121 net121 io_oeb[20] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput143 net143 io_oeb[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput154 net154 io_out[17] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput176 net176 io_out[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput165 net165 io_out[27] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_115_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput187 net187 la_data_out[18] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput198 net198 la_data_out[28] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_116_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input28_I la_data_in[59] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__893__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__657__A1 _203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_884_ net138 net117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput12 la_data_in[43] net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput23 la_data_in[54] net23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput34 la_data_in[65] net34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput45 la_oenb[42] net45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput56 la_oenb[53] net56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput67 la_oenb[64] net67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput78 wbs_dat_i[16] net78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput89 wbs_dat_i[26] net89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__888__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__350__I0 net33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_867_ net138 net109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__653__I1 net150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__644__I1 net177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input95_I wbs_dat_i[31] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_721_ _025_ clknet_3_5__leaf_counter.clk net162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_84_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_652_ _322_ _045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__635__I1 net173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_583_ net26 _263_ _264_ net88 _272_ _273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_16_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_919_ net153 net185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_290 la_data_out[69] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_143_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_3_3__f_counter.clk_I clknet_0_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input10_I la_data_in[41] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_704_ _008_ clknet_3_1__leaf_counter.clk net175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__481__A2 _103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_635_ net238 net173 _309_ _313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_566_ _256_ _257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_497_ _077_ _199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__702__CLK clknet_3_3__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I la_data_in[33] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__472__A2 _173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input58_I la_oenb[55] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__896__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__463__A2 _166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output214_I net214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_420_ _133_ _134_ net71 _076_ _135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__725__CLK clknet_3_4__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_351_ _067_ counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_618_ net66 _151_ _302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_549_ net155 net156 _227_ _242_ _243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_9_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__693__A2 _339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__748__CLK clknet_3_2__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__381__A1 net60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output164_I net164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_403_ net50 _109_ _118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__372__A1 _068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__675__A2 _324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput133 net133 io_oeb[31] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput122 net122 io_oeb[21] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput111 net111 io_oeb[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput166 net166 io_out[28] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput155 net155 io_out[18] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput177 net177 io_out[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput144 net144 io_oeb[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_138_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput188 net188 la_data_out[19] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput199 net199 la_data_out[29] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_29_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__414__I _128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__350__S net67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__657__A2 _324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_883_ net138 net116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput13 la_data_in[44] net13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput35 la_oenb[32] net35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput46 la_oenb[43] net46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput24 la_data_in[55] net24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput68 la_oenb[65] net68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput57 la_oenb[54] net57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput79 wbs_dat_i[17] net79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__584__A1 _246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input40_I la_oenb[37] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__409__I _087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__350__I1 wb_clk_i vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__557__A1 _246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input88_I wbs_dat_i[25] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__899__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_720_ _024_ clknet_3_7__leaf_counter.clk net161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_40_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_651_ net214 net149 _321_ _322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_582_ _265_ _266_ _267_ _271_ _272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_44_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__548__A1 net158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_918_ net152 net184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__539__A1 _231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_280 la_data_out[59] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_291 la_data_out[70] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_132_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__422__I net157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_703_ _007_ clknet_3_3__leaf_counter.clk net174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_634_ _312_ _037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_565_ _142_ _255_ _256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_496_ _172_ _198_ _013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_1__f_counter.clk clknet_0_counter.clk clknet_3_1__leaf_counter.clk vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_131_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_350_ net33 wb_clk_i net67 _067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_617_ _257_ _298_ _300_ _301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_17_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_548_ net158 net159 _242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_479_ _182_ _184_ _185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__390__A2 _101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input105_I wbs_sel_i[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__381__A2 net63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input70_I wbs_cyc_i vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output157_I net157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__436__A3 net96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_402_ net39 net58 _106_ _117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__363__A2 _071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput134 net134 io_oeb[32] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput123 net123 io_oeb[22] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput112 net112 io_oeb[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_12_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput145 net145 io_oeb[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput167 net167 io_out[29] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput156 net156 io_out[19] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_142_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__715__CLK clknet_3_7__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput178 net178 la_data_out[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput189 net189 la_data_out[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_141_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_882_ net138 net115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput36 la_oenb[33] net36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput14 la_data_in[45] net14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput25 la_data_in[56] net25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput69 wb_rst_i net69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput47 la_oenb[44] net47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput58 la_oenb[55] net58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__738__CLK clknet_3_0__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input33_I la_data_in[64] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_934_ net170 net202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__638__I0 net239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__629__I0 net233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__493__A1 net148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_650_ _308_ _321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_72_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_581_ _270_ _271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__548__A2 net159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__484__A1 net147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_917_ net151 net183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__539__A2 net156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_281 la_data_out[60] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_270 la_data_out[49] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_143_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_292 la_data_out[71] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_58_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__466__A1 net108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_702_ _006_ clknet_3_3__leaf_counter.clk net173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_633_ net237 _153_ _309_ _312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_564_ _124_ _254_ _255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_495_ net13 _102_ _175_ _197_ _194_ net74 _198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_32_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_616_ _292_ _294_ _293_ _299_ _300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_17_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_547_ net158 _235_ _241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_17_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_478_ _168_ _169_ _183_ _184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_13_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_counter.clk counter.clk clknet_0_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_141_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__602__A1 net164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__518__I _216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input63_I la_oenb[60] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__436__A4 _138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_401_ _112_ _113_ _114_ _115_ _116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XPHY_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_127_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__596__B1 _279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput124 net124 io_oeb[23] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput113 net113 io_oeb[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_115_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput135 net135 io_oeb[33] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput168 net168 io_out[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput157 net157 io_out[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput146 net146 io_out[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_102_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput179 net179 la_data_out[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_101_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_881_ net138 net114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput37 la_oenb[34] net37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput15 la_data_in[46] net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 la_data_in[57] net26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput48 la_oenb[45] net48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput59 la_oenb[56] net59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__621__I _075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input26_I la_data_in[57] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_933_ net169 net201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__638__I1 net174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__705__CLK clknet_3_6__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__629__I1 net168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__526__I _216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_580_ _247_ _268_ _243_ _269_ _270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__728__CLK clknet_3_7__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_916_ net150 net182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_260 la_data_out[39] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_282 la_data_out[61] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_271 la_data_out[50] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_89_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_293 la_data_out[72] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_144_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input93_I wbs_dat_i[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_701_ _005_ clknet_3_1__leaf_counter.clk net172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_91_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_632_ _311_ _036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_563_ _125_ net106 _254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_494_ net149 _196_ _197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_8_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__384__A1 net48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_615_ net170 _299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_546_ _223_ _240_ _021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_477_ net177 net176 _183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__624__I _074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__602__A2 net165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__366__A1 net59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__534__I net155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input56_I la_oenb[53] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_400_ net41 _070_ _115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__357__A1 _068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__596__A1 net90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_529_ _210_ _203_ _204_ _226_ _227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_92_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__354__I _069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput125 net125 io_oeb[24] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput114 net114 io_oeb[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_133_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput136 net136 io_oeb[34] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput158 net158 io_out[20] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput147 net147 io_out[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_138_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__520__A1 net153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput169 net169 io_out[30] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_115_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__587__A1 _275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output162_I net162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__511__A1 _210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_880_ net138 net113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__439__I _077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput16 la_data_in[47] net16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput27 la_data_in[58] net27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__902__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput38 la_oenb[35] net38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput49 la_oenb[46] net49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__349__I _066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input19_I la_data_in[50] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_932_ net167 net199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_915_ net149 net181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__627__I _074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__362__I _065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_272 la_data_out[51] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_250 irq[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_261 la_data_out[40] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_144_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_283 la_data_out[62] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_294 la_data_out[73] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_143_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input86_I wbs_dat_i[23] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_700_ _004_ clknet_3_3__leaf_counter.clk net171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_631_ net236 net171 _309_ _311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_562_ _246_ _253_ _024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_493_ net148 _192_ _196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_25_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__910__I net175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__393__A2 _106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__718__CLK clknet_3_5__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_614_ net167 net169 net170 _288_ _298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_17_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_545_ net21 _108_ _217_ _239_ _233_ net83 _240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_17_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_476_ net176 _177_ net177 _182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__905__I net168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__686__I0 net230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__602__A3 net166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__523__C1 _221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input49_I la_oenb[46] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__357__A2 _072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__668__I0 net221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_528_ net153 net154 _226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_459_ net175 _167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput115 net115 io_oeb[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_126_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__370__I _069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput137 net137 io_oeb[35] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput126 net126 io_oeb[25] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput159 net159 io_out[21] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput148 net148 io_out[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_86_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input103_I wbs_sel_i[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output155_I net155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput17 la_data_in[48] net17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 la_data_in[59] net28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput39 la_oenb[36] net39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__404__B _109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__569__A2 _254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_931_ net166 net198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__913__I net147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__751__CLK clknet_3_1__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__411__A1 _125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__478__A1 _168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input31_I la_data_in[62] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__402__A1 net39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_914_ net148 net180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__641__A1 _168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__908__I net173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_273 la_data_out[52] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_251 irq[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_262 la_data_out[41] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_32_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_284 la_data_out[63] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_295 la_data_out[74] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__553__I _066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input79_I wbs_dat_i[17] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_630_ _310_ _035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__623__A1 _131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_561_ net24 _250_ _216_ _252_ _233_ net86 _253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_17_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_492_ _172_ _195_ _012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__614__A1 net167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_759_ _063_ clknet_3_3__leaf_counter.clk net234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__605__A1 _274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_613_ _296_ _297_ _188_ _031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_544_ net158 _235_ _239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_17_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_475_ _172_ _181_ _009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__921__I net155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__532__B1 _221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__686__I1 _278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__523__C2 net78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__668__I1 net156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__708__CLK clknet_3_6__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_527_ net153 _218_ net154 _225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__916__I net150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_458_ net42 _165_ _166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_389_ _099_ _100_ _102_ _103_ _104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_13_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput116 net116 io_oeb[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_115_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput138 net138 io_oeb[36] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput127 net127 io_oeb[26] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput149 net149 io_out[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_142_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__347__I0 net34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input61_I la_oenb[58] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output148_I net148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput18 la_data_in[49] net18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput29 la_data_in[60] net29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_930_ net165 net197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__411__A2 net103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__478__A2 _169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input24_I la_data_in[55] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__402__A2 net58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_913_ net147 net179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__641__A2 _000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__924__I net159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_263 la_data_out[42] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_252 irq[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_99_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_285 la_data_out[64] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_274 la_data_out[53] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_296 la_data_out[75] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__396__A1 _105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__623__A2 _000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_560_ net161 _251_ _252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_491_ net12 _092_ _176_ _193_ _194_ net73 _195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_129_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__741__CLK clknet_3_2__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__919__I net153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__614__A2 net169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_758_ _062_ clknet_3_3__leaf_counter.clk net232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__378__A1 net64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_689_ _343_ _061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__550__A1 net159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__369__A1 net62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input91_I wbs_dat_i[28] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output178_I net178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_612_ net31 _095_ _264_ net94 _297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_18_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_543_ _223_ _238_ _020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_474_ net9 _090_ _176_ _178_ _180_ net101 _181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_111_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__532__B2 net79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__532__A1 net18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__599__A1 net166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__523__A1 net17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__514__A1 net51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_526_ _216_ _224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_457_ _072_ _165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_388_ net44 _101_ _103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__932__I net167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__505__B2 _203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput128 net128 io_oeb[27] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput117 net117 io_oeb[17] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput139 net139 io_oeb[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_5_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__347__I1 net69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input54_I la_oenb[51] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output210_I net210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput19 la_data_in[50] net19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__927__I net162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_509_ _199_ _209_ _015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output160_I net160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__420__A3 net71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__482__I _065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__431__B _143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input17_I la_data_in[48] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_912_ net177 net209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_0_counter.clk_I counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_264 la_data_out[43] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_253 la_data_out[32] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_32_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_275 la_data_out[54] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_297 la_data_out[76] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_286 la_data_out[65] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input9_I la_data_in[40] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__396__A2 _107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_1__f_counter.clk_I clknet_0_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__387__A2 _101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_490_ _179_ _194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_757_ _061_ clknet_3_2__leaf_counter.clk net231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__614__A3 net170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_688_ net231 net166 _337_ _343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__369__A2 _071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input84_I wbs_dat_i[21] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_611_ _257_ _291_ _295_ _296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_542_ net20 _091_ _221_ net81 _237_ _238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_2988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_473_ _179_ _180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__532__A2 _112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__599__A2 _279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__665__I _308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__523__A2 _213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__731__CLK clknet_3_0__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__575__I net163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__508__C _208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_108_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__686__S _337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__450__A1 net173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_525_ _066_ _223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_456_ _150_ _164_ _007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_387_ net47 _101_ _102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__754__CLK clknet_3_3__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput129 net129 io_oeb[28] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput118 net118 io_oeb[18] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_141_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_6__f_counter.clk_I clknet_0_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__441__A1 net39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input47_I la_oenb[44] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output203_I net203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__499__A1 net150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__423__A1 _136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_508_ net76 _180_ _205_ _206_ _208_ _209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_92_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_439_ _077_ _150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input101_I wbs_dat_i[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output153_I net153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__420__A4 _076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__571__C2 net87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_911_ net176 net208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_243 io_oeb[37] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_116_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_254 la_data_out[33] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_265 la_data_out[44] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_276 la_data_out[55] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_287 la_data_out[66] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_143_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_298 la_data_out[77] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_98_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__396__A3 _108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__608__A1 _275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__578__I net161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__631__I1 net171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__527__B net154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_756_ _060_ clknet_3_6__leaf_counter.clk net230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__614__A4 _288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_687_ _342_ _060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input77_I wbs_dat_i[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output233_I net233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_610_ _292_ _293_ _294_ _295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_541_ _224_ _235_ _236_ _237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_17_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_472_ _156_ _173_ _179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_739_ _043_ clknet_3_0__leaf_counter.clk net212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__681__I _076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__540__B net156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_524_ _199_ _222_ _017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_455_ net7 _115_ _128_ _163_ _157_ net99 _164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_144_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_386_ _085_ _101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput119 net119 io_oeb[19] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_142_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_3_4__f_counter.clk clknet_0_counter.clk clknet_3_4__leaf_counter.clk vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_20_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__586__I net164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__423__A2 _130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_507_ net49 _207_ _165_ _208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_14_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__721__CLK clknet_3_5__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_438_ net138 _149_ _004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_369_ net62 _071_ _083_ _084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output146_I net146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__405__A2 net51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__744__CLK clknet_3_0__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__580__A1 _247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__571__A1 net25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_910_ net175 net207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__562__A1 _246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_example_244 io_out[32] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_128_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_255 la_data_out[34] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_99_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_266 la_data_out[45] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_277 la_data_out[56] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_288 la_data_out[67] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_299 la_data_out[78] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__396__A4 _110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__608__A2 _278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input22_I la_data_in[53] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__544__A1 net158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_755_ _059_ clknet_3_2__leaf_counter.clk net229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_686_ net230 _278_ _337_ _342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__437__C _148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__535__A1 _231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_540_ _231_ _228_ net156 _236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_471_ net176 _177_ _178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_13_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_738_ _042_ clknet_3_0__leaf_counter.clk net242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_669_ _332_ _052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__508__A1 net76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__872__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output176_I net176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_523_ net17 _213_ _217_ _219_ _221_ net78 _222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_144_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_454_ net174 _162_ _163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_2798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_385_ net45 _086_ _100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput109 net109 io_oeb[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_115_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__426__B1 _129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__867__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__417__B1 _129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__432__A3 net93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_506_ net15 _207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_437_ net4 _113_ _129_ _147_ _148_ _149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_14_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_368_ _081_ _082_ _083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__696__CLK clknet_3_1__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input52_I la_oenb[49] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__580__A2 _268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__399__A2 _109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_64_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__880__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__711__CLK clknet_3_7__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_245 io_out[33] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_144_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_267 la_data_out[46] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_278 la_data_out[57] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_256 la_data_out[35] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_289 la_data_out[68] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_97_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__625__I0 net222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__734__CLK clknet_3_1__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__608__A3 net166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__875__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input15_I la_data_in[46] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_754_ _058_ clknet_3_3__leaf_counter.clk net228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_685_ _341_ _059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__757__CLK clknet_3_2__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input7_I la_data_in[38] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__471__A1 net176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__462__A1 _168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output219_I net219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_470_ _168_ _169_ _177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__453__A1 net173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_737_ _041_ clknet_3_2__leaf_counter.clk net241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_668_ net221 net156 _330_ _332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_599_ net166 _279_ _286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_32_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__444__A1 _153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input82_I wbs_dat_i[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output169_I net169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__683__A1 _265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__435__A1 net171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_522_ _220_ _221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_453_ net173 _153_ _154_ _162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_14_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_384_ net48 _086_ _099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__674__A1 net225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__426__A1 net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__417__B2 _131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__417__A1 net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__432__A4 _138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__883__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_505_ _142_ _174_ _204_ _203_ _206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_436_ _133_ _134_ net96 _138_ _148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_13_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_367_ net37 _080_ _082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__647__A1 _191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__670__I1 net158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__878__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input45_I la_oenb[42] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_3_0__f_counter.clk clknet_0_counter.clk clknet_3_0__leaf_counter.clk vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__661__I1 net153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_419_ net103 _134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__556__C2 net85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__556__B1 _216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output151_I net151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_246 io_out[34] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_11_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_268 la_data_out[47] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_279 la_data_out[58] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_257 la_data_out[36] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_899_ net138 net134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__625__I1 _136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__891__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_753_ _057_ clknet_3_6__leaf_counter.clk net227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_684_ net229 _275_ _337_ _341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__701__CLK clknet_3_1__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__886__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__462__A2 _169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__453__A2 _153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_736_ _040_ clknet_3_0__leaf_counter.clk net240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_667_ _331_ _051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_598_ net63 _151_ _285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__724__CLK clknet_3_5__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__692__A2 _306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__380__A1 net65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input75_I wbs_dat_i[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__683__A2 _339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output231_I net231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__435__A2 _141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__747__CLK clknet_3_2__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_521_ _156_ _214_ _220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_452_ _150_ _161_ _006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_383_ _090_ _091_ _092_ _097_ _098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_144_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__674__A2 _326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__426__A2 _088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_719_ _023_ clknet_3_7__leaf_counter.clk net160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__417__A2 _078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__656__A2 _304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_504_ _203_ _204_ _205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_33_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_435_ net171 _141_ _147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_13_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_366_ net59 _080_ _081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__592__A1 _275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__647__A2 _000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__583__B2 net88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__583__A1 net26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input38_I la_oenb[35] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__894__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_418_ _125_ _133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_349_ _066_ net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_128_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__556__A1 net23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__889__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__547__A1 net158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_247 io_out[35] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_258 la_data_out[37] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_269 la_data_out[48] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_32_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_898_ net138 net133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__483__B _188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__502__I net151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__474__C2 net101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__529__A1 _210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_752_ _056_ clknet_3_1__leaf_counter.clk net226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_683_ _265_ _339_ _340_ _058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__447__C2 net97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__447__B1 _129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input20_I la_data_in[51] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_735_ _039_ clknet_3_2__leaf_counter.clk net239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_666_ net220 _231_ _330_ _331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_597_ _274_ _284_ _028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__699__CLK clknet_3_3__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input68_I la_oenb[65] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__897__I net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_520_ net153 _218_ _219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_6_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output224_I net224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_451_ net6 _110_ _128_ _160_ _157_ net98 _161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_26_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_382_ _093_ _094_ _095_ _096_ _097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_13_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_718_ _022_ clknet_3_5__leaf_counter.clk net159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_649_ _320_ _044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__510__I net152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output174_I net174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__714__CLK clknet_3_4__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_503_ net150 net149 net148 _192_ _204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_2587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_434_ net138 _146_ _003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_365_ _079_ _080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__737__CLK clknet_3_2__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__415__I net146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_417_ net1 _078_ _129_ _131_ _132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_15_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_348_ _065_ _066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__556__A2 _107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input50_I la_oenb[47] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput240 net240 wbs_dat_o[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_248 io_out[36] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_259 la_data_out[38] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_136_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_897_ net138 net132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__474__A1 net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__529__A2 _203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input98_I wbs_dat_i[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_751_ _055_ clknet_3_1__leaf_counter.clk net225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_682_ net228 _326_ _340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__695__A1 _299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__447__A1 net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input13_I la_data_in[44] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__438__A1 net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_734_ _038_ clknet_3_1__leaf_counter.clk net238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_665_ _308_ _330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_16_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_596_ net90 _264_ _279_ _281_ _283_ _284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__610__A1 _292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__677__A1 _268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I la_data_in[36] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__601__A1 _274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_450_ net173 _159_ _160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__418__I _125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_381_ net60 net63 _070_ _096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_717_ _021_ clknet_3_4__leaf_counter.clk net158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_17_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_648_ net213 net148 _314_ _320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_579_ net162 net163 _269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input80_I wbs_dat_i[18] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output167_I net167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_502_ net151 _203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_2588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_433_ net3 _082_ _141_ _144_ _145_ _146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_26_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__592__B _278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_364_ _069_ _079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_416_ _130_ _131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_347_ net34 net69 net68 _065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__704__CLK clknet_3_1__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput241 net241 wbs_dat_o[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput230 net230 wbs_dat_o[27] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input43_I la_oenb[40] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_249 io_out[37] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_109_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_896_ net138 net130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__727__CLK clknet_3_7__leaf_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__474__A2 _090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_750_ _054_ clknet_3_2__leaf_counter.clk net224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_681_ _076_ _339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_879_ net138 net112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__695__A2 _339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__447__A2 _152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__383__A1 _090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_733_ _037_ clknet_3_1__leaf_counter.clk net237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_664_ _329_ _050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_595_ net62 _282_ _072_ _283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_32_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__374__A1 _087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__677__A2 _324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_380_ net65 _079_ _095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__659__A2 _326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_716_ _020_ clknet_3_4__leaf_counter.clk net156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_131_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__609__I net169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_647_ _191_ _000_ _319_ _043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__595__A1 net62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_578_ net161 _268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_3_4__f_counter.clk_I clknet_0_counter.clk vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

