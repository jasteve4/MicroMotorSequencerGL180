* NGSPICE file created from controller_core.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

.subckt controller_core clock clock_out[0] clock_out[1] clock_out[2] clock_out[3]
+ clock_out[4] clock_out[5] clock_out[6] clock_out[7] clock_out[8] clock_out[9] col_select_left[0]
+ col_select_left[1] col_select_left[2] col_select_left[3] col_select_left[4] col_select_left[5]
+ col_select_right[0] col_select_right[1] col_select_right[2] col_select_right[3]
+ col_select_right[4] col_select_right[5] data_out_left[0] data_out_left[10] data_out_left[11]
+ data_out_left[12] data_out_left[13] data_out_left[14] data_out_left[15] data_out_left[1]
+ data_out_left[2] data_out_left[3] data_out_left[4] data_out_left[5] data_out_left[6]
+ data_out_left[7] data_out_left[8] data_out_left[9] data_out_right[0] data_out_right[10]
+ data_out_right[11] data_out_right[12] data_out_right[13] data_out_right[14] data_out_right[15]
+ data_out_right[1] data_out_right[2] data_out_right[3] data_out_right[4] data_out_right[5]
+ data_out_right[6] data_out_right[7] data_out_right[8] data_out_right[9] inverter_select[0]
+ inverter_select[1] inverter_select[2] inverter_select[3] inverter_select[4] inverter_select[5]
+ inverter_select[6] inverter_select[7] inverter_select[8] inverter_select[9] io_control_trigger_in
+ io_control_trigger_oeb io_driver_io_oeb[0] io_driver_io_oeb[10] io_driver_io_oeb[11]
+ io_driver_io_oeb[12] io_driver_io_oeb[13] io_driver_io_oeb[14] io_driver_io_oeb[15]
+ io_driver_io_oeb[16] io_driver_io_oeb[17] io_driver_io_oeb[18] io_driver_io_oeb[19]
+ io_driver_io_oeb[1] io_driver_io_oeb[2] io_driver_io_oeb[3] io_driver_io_oeb[4]
+ io_driver_io_oeb[5] io_driver_io_oeb[6] io_driver_io_oeb[7] io_driver_io_oeb[8]
+ io_driver_io_oeb[9] io_latch_data_in io_latch_data_oeb io_reset_n_in io_reset_n_oeb
+ io_update_cycle_complete_oeb io_update_cycle_complete_out la_data_in[0] la_data_in[10]
+ la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[1] la_data_in[2] la_data_in[3] la_data_in[4] la_data_in[5]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_oenb[0] la_oenb[10] la_oenb[11]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[1]
+ la_oenb[2] la_oenb[3] la_oenb[4] la_oenb[5] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9]
+ mem_address_left[0] mem_address_left[1] mem_address_left[2] mem_address_left[3]
+ mem_address_left[4] mem_address_left[5] mem_address_left[6] mem_address_left[7]
+ mem_address_left[8] mem_address_left[9] mem_address_right[0] mem_address_right[1]
+ mem_address_right[2] mem_address_right[3] mem_address_right[4] mem_address_right[5]
+ mem_address_right[6] mem_address_right[7] mem_address_right[8] mem_address_right[9]
+ mem_write_n[0] mem_write_n[1] mem_write_n[2] mem_write_n[3] mem_write_n[4] mem_write_n[5]
+ mem_write_n[6] mem_write_n[7] mem_write_n[8] mem_write_n[9] output_active_left output_active_right
+ row_col_select[0] row_col_select[1] row_col_select[2] row_col_select[3] row_col_select[4]
+ row_col_select[5] row_col_select[6] row_col_select[7] row_col_select[8] row_col_select[9]
+ row_select_left[0] row_select_left[1] row_select_left[2] row_select_left[3] row_select_left[4]
+ row_select_left[5] row_select_right[0] row_select_right[1] row_select_right[2] row_select_right[3]
+ row_select_right[4] row_select_right[5] spi_data[0] spi_data[10] spi_data[11] spi_data[12]
+ spi_data[13] spi_data[14] spi_data[15] spi_data[16] spi_data[17] spi_data[18] spi_data[19]
+ spi_data[1] spi_data[20] spi_data[21] spi_data[22] spi_data[23] spi_data[24] spi_data[25]
+ spi_data[26] spi_data[27] spi_data[28] spi_data[29] spi_data[2] spi_data[30] spi_data[31]
+ spi_data[3] spi_data[4] spi_data[5] spi_data[6] spi_data[7] spi_data[8] spi_data[9]
+ spi_data_clock vccd1 vssd1
XTAP_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3155_ spi_data_crossing\[18\].A clknet_leaf_8_clock spi_data_crossing\[18\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3086_ _0220_ clknet_leaf_5_clock u1.timer\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2106_ _0402_ _0493_ _0495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2037_ u1.ccr1\[31\] _0389_ _0426_ _0446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2403__B1 _0691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2939_ _0081_ clknet_leaf_34_clock u1.ordering_complete\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1757__A2 _1342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2706__A1 _0958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3132__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3171__D spi_data_crossing\[26\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1996__A2 _0394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2796__I1 _0363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1942__I u0.cmd\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2712__A4 _0961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2476__A3 _1085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2773__I net8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2722__B _0282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3005__CLK clknet_leaf_35_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2724_ _0968_ _0973_ _0974_ _0237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2655_ u1.ccr1\[18\] _0920_ _0921_ _0922_ _0923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_8_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1606_ _1223_ _1224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3155__CLK clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2586_ _1153_ _0864_ _0865_ spi_data_crossing\[29\].data_sync _0867_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2164__A2 _0530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1537_ _1157_ u0.latch_cmd vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1911__A2 _0361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1468_ _1072_ _1093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3207_ _0277_ clknet_leaf_38_clock net159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3138_ net41 net72 spi_data_crossing\[10\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2683__I _0933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3069_ _0210_ clknet_leaf_13_clock u1.row_sel\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1969__A2 _0400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3028__CLK clknet_leaf_31_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2091__A1 u0.cmd\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3178__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2440_ _0754_ _0755_ _0734_ _0759_ _0760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1672__I u1.timer\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2371_ _1100_ _0694_ _0699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_42_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1657__A1 _1247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2707_ _1311_ _0961_ _0963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2638_ u1.ccr1\[11\] _1269_ u1.ccr1\[10\] _1268_ _0906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2569_ _0856_ _0200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1582__I u1.ccr1\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input36_I la_oenb[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3302__I net168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2128__A2 _0500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_15_clock_I clknet_2_1__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2300__A2 _0627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1940_ u0.cmd\[12\] _0383_ _0384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1871_ u1.col_sel\[0\] _0332_ _0334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2423_ u1.ordering_timer\[20\] _0719_ _0734_ _0744_ _0745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2354_ _1103_ _0683_ _0684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2285_ u1.ordering_timer\[4\] _0623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1802__A1 _0281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2358__A2 _0687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2201__I _0552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1869__A1 _1212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2294__A1 _0611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1487__I u1.ordering_complete\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2860__CLK clknet_leaf_7_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3216__CLK clknet_leaf_22_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2070_ _0471_ _0086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2972_ _0114_ clknet_leaf_14_clock u1.row_limit\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2588__A2 _0864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1923_ u0.cmd\[7\] _0372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_19_clock clknet_2_3__leaf_clock clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1854_ u1.col_sel\[1\] _0317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1785_ u0.timer_enable _1402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2406_ _0729_ _0723_ _0730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2337_ _0669_ _0155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2268_ _0599_ _0601_ _0604_ _0608_ _0609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2199_ _0551_ _0135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2028__A1 _0381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2883__CLK clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3239__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2640__B _0907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2200__A1 u0.cmd\[19\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2019__A1 _0372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1490__A2 _1110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1778__B1 _1344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1945__I u0.cmd\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1570_ u1.timer\[6\] _1188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3240_ u0.cmd\[22\] clknet_leaf_10_clock net168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3171_ spi_data_crossing\[26\].A clknet_leaf_10_clock spi_data_crossing\[26\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2122_ u1.ordering_complete\[26\] _0504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2053_ _0399_ _0459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2217__S _0558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1481__A2 u1.ordering_complete\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2955_ _0097_ clknet_leaf_33_clock u1.ordering_complete\[17\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2886_ _0020_ clknet_leaf_12_clock u0.mem_write_n\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1906_ u0.cmd\[2\] _0360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1837_ _0302_ _0303_ _0305_ _0018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2033__I1 _0385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2733__A2 _0978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1768_ _1256_ u1.ccr0\[15\] _1306_ _1385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1699_ _1302_ _1308_ _1309_ _1315_ _1316_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2497__A1 _1082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output105_I net105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3310__I net207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3061__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3169__D spi_data_crossing\[25\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2421__A1 u1.ordering_complete\[20\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2024__I1 _0376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput75 net75 clock_out[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput86 net86 col_select_left[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_49_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput97 net97 data_out_left[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_48_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2037__S _0426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2660__A1 u1.ccr1\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2740_ _0983_ _0984_ _0985_ _0242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2671_ _0933_ _0937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1622_ u1.ccr1\[18\] u1.timer\[18\] _1240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2015__I1 _0367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1518__A3 _1137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1553_ u1.timer\[31\] _1171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1484_ u1.ordering_timer\[9\] _1109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3223_ u1.inverter_select\[9\] clknet_leaf_22_clock net136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3154_ net49 net72 spi_data_crossing\[18\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3085_ _0219_ clknet_leaf_38_clock net149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2105_ _1067_ _0489_ _0494_ _0098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2036_ _0445_ _0078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3084__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2651__A1 _1227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2403__A1 _1068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2938_ _0080_ clknet_leaf_34_clock u1.ordering_complete\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2869_ _0026_ clknet_leaf_18_clock u1.col_sel\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2921__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2006__I1 _0360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input66_I spi_data[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2706__A2 _0961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1534__B _1155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3305__I net171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2190__I0 _0367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_2_1__f_clock_I clknet_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2181__I0 _0517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2476__A4 _0784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2944__CLK clknet_leaf_2_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2723_ _0282_ u1.timer\[16\] _0970_ _0974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2654_ _0429_ u1.timer\[19\] _0922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2585_ _0866_ _0206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1605_ u1.timer\[20\] _1223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1536_ _1156_ u0.u11.impulse_gen\[1\] _1157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1467_ _1088_ u1.ordering_complete\[25\] _1091_ _1092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_28_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3206_ _0276_ clknet_leaf_27_clock u1.ccr0\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3137_ spi_data_crossing\[9\].A clknet_leaf_2_clock spi_data_crossing\[9\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3068_ _0023_ clknet_leaf_7_clock u1.output_active vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2624__A1 _0890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2019_ _0372_ _0431_ _0436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3182__D _0252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2615__A1 u1.row_sel\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1418__A2 u0.cmd\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2967__CLK clknet_leaf_33_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2091__A2 _0478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_11_clock_I clknet_2_1__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2370_ u1.ordering_timer\[14\] _0698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2082__A2 _0453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3122__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2706_ _0958_ _0961_ _0962_ _0231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xoutput210 net210 row_select_right[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2637_ _0905_ net38 _0219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2568_ u0.cmd\[22\] _0852_ _0853_ spi_data_crossing\[22\].data_sync _0856_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1896__A2 _0348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1519_ _1070_ _1095_ _1120_ _1143_ _1144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_2499_ u1.ordering_timer\[31\] _0810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2145__I0 _0459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input29_I la_oenb[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3177__D spi_data_crossing\[29\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output97_I net97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3145__CLK clknet_leaf_2_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1948__I u0.cmd\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1870_ u1.col_sel\[0\] _0332_ _0333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1683__I u1.timer\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2422_ _0735_ _0742_ _0743_ _0744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2353_ _0675_ _0677_ _0683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2284_ _0622_ _0149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1802__A2 _1322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1999_ _0422_ _0423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_14_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1566__B2 _1165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1566__A1 u1.ccr1\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3018__CLK clknet_leaf_35_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1869__A2 _0309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2118__I0 _0474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2818__A1 u0.cmd\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3168__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2109__I0 _0464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2971_ _0113_ clknet_leaf_14_clock u1.row_limit\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1922_ _1329_ _0359_ _0371_ _0038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1853_ u1.col_sel\[2\] _0316_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1784_ _1292_ _1374_ _1400_ _1401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2405_ _1065_ _0729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2336_ u1.ordering_timer\[9\] _0655_ _0662_ _0668_ _0669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2267_ u1.ordering_complete\[1\] _0605_ _0607_ _0608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2198_ _0476_ u1.inverter_select\[9\] _0539_ _0551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2276__A2 _0597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2028__A2 _0423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3190__D _0260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2019__A2 _0431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1778__A1 _1394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1778__B2 _1345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2122__I u1.ordering_complete\[26\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1950__A1 _1352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1961__I u0.cmd\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3170_ net58 net72 spi_data_crossing\[26\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2121_ _0503_ _0105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2052_ _1134_ _0453_ _0458_ _0081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2954_ _0096_ clknet_leaf_34_clock u1.ordering_complete\[16\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2885_ _0019_ clknet_leaf_11_clock u0.mem_write_n\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1905_ _0358_ _0359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1836_ _0301_ _0305_ _0017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1767_ _1302_ _1308_ _1384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1698_ _1312_ _1314_ _1315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2497__A2 _0716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2319_ _0653_ _0153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3299_ net165 net175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2850__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input11_I la_data_in[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3206__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2421__A2 _0687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3185__D _0255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2724__A3 _0974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput76 net76 clock_out[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput98 net98 data_out_left[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput87 net87 col_select_left[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__2488__A2 _0796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_18_clock clknet_2_3__leaf_clock clknet_leaf_18_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2670_ _0935_ _0936_ _0221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1621_ u1.ccr1\[19\] u1.timer\[19\] _1239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_8_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1552_ u1.ccr1\[25\] _1164_ u1.ccr1\[24\] _1166_ _1169_ _1170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__2787__I _1013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1483_ _1099_ _1102_ _1107_ _1108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3222_ u1.inverter_select\[8\] clknet_leaf_21_clock net135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2873__CLK clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3153_ spi_data_crossing\[17\].A clknet_leaf_8_clock spi_data_crossing\[17\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input3_I io_reset_n_in vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2479__A2 _0711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2104_ _0399_ _0493_ _0494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3084_ _0010_ clknet_leaf_9_clock u0.run_state\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3229__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2035_ u1.ccr1\[30\] _0387_ _0438_ _0445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2100__A1 _1060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2403__A2 _0719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2937_ _0079_ clknet_leaf_27_clock u1.ccr1\[31\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1866__I _1402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2868_ _0025_ clknet_leaf_18_clock u1.col_sel\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1819_ u0.cmd\[30\] _0295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2167__A1 _0399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2799_ _0404_ _1021_ _1022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input59_I spi_data[27] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output215_I net215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2896__CLK clknet_leaf_25_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2633__A2 latch_data vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1686__I u1.timer\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2722_ _0283_ _0971_ _0282_ _0973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2397__A1 _1068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2653_ _1241_ _1238_ _1242_ _0921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2584_ u0.cmd\[28\] _0864_ _0865_ spi_data_crossing\[28\].data_sync _0866_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1604_ _1202_ _1211_ _1221_ _1222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_12_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1535_ u0.u11.impulse_gen\[0\] _1156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1466_ u1.ordering_timer\[24\] _1086_ _1091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3205_ _0275_ clknet_leaf_27_clock u1.ccr0\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3051__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3136_ net71 net72 spi_data_crossing\[9\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3067_ _0209_ clknet_leaf_9_clock u0.cmd\[31\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2018_ _1226_ _0430_ _0435_ _0070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output165_I net165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2560__B2 spi_data_crossing\[19\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2560__A1 u0.cmd\[19\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2615__A2 _0875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1418__A3 _1042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3074__CLK clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2911__CLK clknet_leaf_7_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2705_ _1272_ _0959_ _0962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput200 net200 row_col_select[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2636_ net20 _0905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput211 net211 row_select_right[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2567_ _0855_ _0199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2542__A1 _0442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1518_ _1132_ _1135_ _1137_ _1142_ _1143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_2498_ _0565_ _0601_ _0808_ _0809_ _0176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2542__B2 spi_data_crossing\[12\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1449_ u1.ordering_timer\[31\] _1073_ _1074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2145__I1 u1.row_limit\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3119_ spi_data_crossing\[0\].A clknet_leaf_38_clock spi_data_crossing\[0\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3097__CLK clknet_leaf_4_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2934__CLK clknet_leaf_28_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2125__I u1.ordering_complete\[27\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2072__I0 _0472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2061__S _0460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2421_ u1.ordering_complete\[20\] _0687_ _0743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2524__A1 _0466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2352_ _0625_ _0682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2524__B2 spi_data_crossing\[5\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2283_ u1.ordering_timer\[3\] _0601_ _0604_ _0621_ _0622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1802__A3 _0282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1998_ _0346_ _0391_ _0351_ _0422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__2763__A1 _1351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1566__A2 _1173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2619_ u1.row_sel\[2\] u1.row_sel\[1\] _0892_ _0895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2957__CLK clknet_leaf_33_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input41_I spi_data[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2118__I1 u1.ordering_complete\[24\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2818__A2 _1029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output128_I net128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3188__D _0258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1985__S _0397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2109__I1 u1.ordering_complete\[20\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3112__CLK clknet_leaf_24_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1493__A1 _1111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1959__I _0393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2970_ _0112_ clknet_leaf_14_clock u1.row_limit\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1921_ _0369_ _0370_ _0371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1852_ _0313_ u1.col_limit\[3\] _0314_ u1.col_limit\[4\] _0315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_30_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1783_ _1362_ _1393_ _1399_ _1400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2745__A1 _0983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2404_ _0728_ _0163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2335_ _0643_ _0666_ _0667_ _0668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2266_ _0606_ _0607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2197_ _0550_ _0134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3135__CLK clknet_leaf_2_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2727__A1 _0968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1950__A2 _0361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2120_ _0476_ u1.ordering_complete\[25\] _0488_ _0503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2051_ _0457_ _0455_ _0458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2953_ _0095_ clknet_leaf_35_clock u1.ordering_complete\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1904_ _0352_ _0358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3008__CLK clknet_leaf_1_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2884_ _0018_ clknet_leaf_11_clock u0.mem_write_n\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1835_ _0298_ _0305_ _0016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3158__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1766_ _1313_ _1382_ _1312_ _1383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1697_ _1267_ u1.ccr0\[8\] _1313_ _1314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1941__A2 _0378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2318_ _0648_ _0626_ _0635_ _0652_ _0653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3298_ net164 net174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2249_ _1080_ _0591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2223__I _1402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2709__A1 _0958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput99 net99 data_out_left[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput77 net77 clock_out[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput88 net88 col_select_left[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2488__A3 _1093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1620__B2 _1237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1620_ u1.ccr1\[17\] _1236_ u1.ccr1\[16\] _1237_ _1238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2176__A2 _0530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1972__I _0393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1551_ u1.ccr1\[30\] _1167_ u1.ccr1\[29\] _1168_ _1169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1482_ _1103_ u1.ordering_complete\[12\] _1105_ _1106_ _1107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3221_ u1.inverter_select\[7\] clknet_leaf_21_clock net134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3152_ net48 net72 spi_data_crossing\[17\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2103_ _0487_ _0493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3083_ _0009_ clknet_leaf_12_clock u0.run_state\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2736__C _0982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2034_ _0444_ _0077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2100__A2 _0489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2936_ _0078_ clknet_leaf_28_clock u1.ccr1\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2867_ _0024_ clknet_leaf_38_clock net160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1818_ _0294_ _0005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2798_ _1011_ _1021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1749_ _1363_ u1.ccr0\[1\] _1365_ _1366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output110_I net110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2064__S _0460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2721_ _1279_ _0932_ _0971_ _0283_ _0972_ _0236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2397__A2 _1059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2652_ _0429_ _1318_ _1321_ _0920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2840__CLK clknet_leaf_18_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2583_ _0846_ _0865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1603_ _1212_ _1216_ _1217_ _1220_ _1221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1534_ _1153_ _1154_ _1155_ _0006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2990__CLK clknet_leaf_22_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3204_ _0274_ clknet_leaf_16_clock u1.ccr0\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1465_ _1085_ _1086_ _1089_ _1090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3135_ spi_data_crossing\[8\].A clknet_leaf_2_clock spi_data_crossing\[8\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3066_ _0208_ clknet_leaf_9_clock u0.cmd\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2017_ _0369_ _0431_ _0435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1832__A1 _0299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2919_ _0061_ clknet_leaf_34_clock u1.ccr1\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_17_clock clknet_2_3__leaf_clock clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input71_I spi_data[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2863__CLK clknet_leaf_15_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3219__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2411__I _0634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2303__A2 _0630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2704_ _1272_ u1.timer\[10\] _0950_ _0955_ _0961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
Xoutput201 net201 row_col_select[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__2790__A2 _1014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2635_ _1156_ _0815_ _0218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput212 net212 row_select_right[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__2321__I _0625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2566_ u0.cmd\[21\] _0852_ _0853_ spi_data_crossing\[21\].data_sync _0855_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2497_ _1082_ _0716_ _0809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1517_ _1139_ u1.ordering_complete\[0\] _1140_ _1141_ _1142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1448_ u1.ordering_complete\[31\] _1073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3118_ net40 net72 spi_data_crossing\[0\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3049_ _0191_ clknet_leaf_3_clock u0.cmd\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2886__CLK clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3041__CLK clknet_leaf_7_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2420_ _1050_ _0737_ _0742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3191__CLK clknet_leaf_16_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2351_ _0681_ _0157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2282_ _0611_ _0619_ _0620_ _0621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1802__A4 _0283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1997_ _1252_ _0400_ _0421_ _0063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2618_ _0891_ _0894_ _0211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1890__I u0.cmd\[16\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2549_ _0843_ _0193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input34_I la_oenb[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3064__CLK clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2901__CLK clknet_leaf_29_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2506__A2 u0.latch_cmd vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1493__A2 _1112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1920_ _0353_ _0370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1851_ u1.col_sel\[4\] _0314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1975__I _0397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2072__S _0470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1782_ _1171_ u1.ccr0\[31\] _1354_ _1398_ _1399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2403_ _1068_ _0719_ _0691_ _0727_ _0728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2334_ _1110_ _0658_ _0667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2265_ _0596_ _0606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2196_ _0474_ u1.inverter_select\[8\] _0539_ _0550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3087__CLK clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2046__I u0.cmd\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2808__I0 u1.ccr0\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2490__B _0709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1641__C1 u1.ccr1\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2924__CLK clknet_leaf_26_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2672__A1 _1364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2360__B1 _0662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2050_ u0.cmd\[1\] _0457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2663__B2 _0930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2947__CLK clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2952_ _0094_ clknet_leaf_35_clock u1.ordering_complete\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1903_ _0357_ _0033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2883_ _0017_ clknet_leaf_13_clock u0.mem_write_n\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1834_ _0304_ u0.cmd\[29\] _0305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1765_ _1294_ _1297_ _1299_ _1309_ _1382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1696_ _1262_ _1310_ _1313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3297_ net163 net173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2317_ _0643_ _0650_ _0651_ _0652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2248_ _1084_ _0589_ _0590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2485__B _0603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2179_ _0513_ u1.inverter_select\[0\] _0540_ _0541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2654__A1 _0429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2406__A1 _0729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3102__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2709__A2 _0963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2590__B1 _0865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3252__CLK clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput89 net89 col_select_right[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput78 net78 clock_out[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1696__A2 _1310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2342__B1 _0662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1620__A2 _1236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1550_ u1.timer\[29\] _1168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1481_ _1101_ u1.ordering_complete\[13\] _1103_ u1.ordering_complete\[12\] _1106_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3220_ u1.inverter_select\[6\] clknet_leaf_21_clock net133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3151_ spi_data_crossing\[16\].A clknet_leaf_7_clock spi_data_crossing\[16\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2102_ _1061_ _0489_ _0492_ _0097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3082_ _0008_ clknet_leaf_9_clock u0.run_state\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2033_ u1.ccr1\[29\] _0385_ _0438_ _0444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3125__CLK clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2935_ _0077_ clknet_leaf_28_clock u1.ccr1\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2866_ reset_n_sync\[0\] clknet_leaf_37_clock reset_n_sync\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2324__I _0629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1817_ u0.cmd\[29\] u0.run_state\[0\] _1155_ _0294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2797_ _1020_ _0264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1748_ _1363_ u1.ccr0\[1\] u1.ccr0\[0\] _1364_ _1365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1679_ u1.ccr0\[10\] _1296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2627__A1 _0890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output103_I net103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2618__A1 _0891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3148__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2633__A4 _1042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2720_ _0283_ _0971_ _0972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2651_ _1227_ _1231_ _0919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1602_ _1218_ _1219_ _1220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2582_ _0844_ _0864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1533_ _1040_ u0.cmd\[30\] _1042_ _1155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_5_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1464_ _1087_ u1.ordering_complete\[26\] _1088_ u1.ordering_complete\[25\] _1089_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3203_ _0273_ clknet_leaf_7_clock u1.ccr0\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_0_clock clock clknet_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3134_ net70 net72 spi_data_crossing\[8\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3065_ _0207_ clknet_leaf_12_clock u0.cmd\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2016_ _0434_ _0069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1832__A2 _1160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2918_ _0060_ clknet_leaf_34_clock u1.ccr1\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2849_ u0.cmd\[5\] clknet_leaf_20_clock net106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1893__I u0.cmd\[19\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input64_I spi_data[31] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2229__I _1096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2139__I _0514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2075__S _0470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2703_ _0958_ _0959_ _0960_ _0230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2634_ _0904_ _0217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput213 net213 row_select_right[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput202 net202 row_col_select[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_47_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2565_ _0854_ _0198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1516_ _1136_ u1.ordering_complete\[2\] _1141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2496_ _0804_ _0807_ _0808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1447_ u1.ordering_timer\[27\] _1072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3117_ _0251_ clknet_leaf_29_clock u1.timer\[31\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3048_ _0190_ clknet_leaf_3_clock u0.cmd\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_2_0__f_clock_I clknet_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output170_I net170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2049__A2 _0453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2980__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1980__A1 u0.cmd\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2350_ _0675_ _0655_ _0662_ _0680_ _0681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_2_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2281_ u1.ordering_complete\[3\] _0597_ _0620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_16_clock clknet_2_2__leaf_clock clknet_leaf_16_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_21_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1996_ _0389_ _0394_ _0421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2617_ _0878_ _0892_ _0894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2548_ _0389_ _0838_ _0839_ spi_data_crossing\[15\].data_sync _0843_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2479_ _0506_ _0711_ _0794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2853__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input27_I la_oenb[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3209__CLK clknet_leaf_38_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output95_I net95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1714__A1 _1327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1850_ u1.col_sel\[3\] _0313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1781_ _1360_ _1397_ _1398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2402_ _1061_ _0720_ _0726_ _0727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2876__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2333_ _0664_ _0665_ _0666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2264_ _1138_ _0599_ _0605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2195_ _0549_ _0133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2681__A2 _0942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2808__I1 _0374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1979_ _1199_ _0409_ _0411_ _0055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3031__CLK clknet_leaf_30_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2672__A2 _1363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3181__CLK clknet_leaf_10_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2173__S _0529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2727__A3 _0976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2899__CLK clknet_leaf_26_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1935__A1 _1344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2700__I _0945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2415__A2 _0737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2951_ _0093_ clknet_leaf_3_clock u1.ordering_complete\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1902_ u1.ccr0\[17\] _0356_ _0354_ _0357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2882_ _0016_ clknet_leaf_13_clock u0.mem_write_n\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1833_ u0.cmd\[28\] _0304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1764_ _1377_ _1378_ _1380_ _1381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1695_ _1300_ _1301_ _1310_ _1311_ _1312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3054__CLK clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3296_ net162 net172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2316_ u1.ordering_complete\[7\] _0630_ _0651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2247_ u1.ordering_timer\[27\] _0506_ u1.ordering_timer\[26\] _0504_ _1089_ _1092_
+ _0589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_22_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2178_ _0539_ _0540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2654__A2 u1.timer\[19\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2057__I _0402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2406__A2 _0723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2590__B2 spi_data_crossing\[31\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2520__I _0817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput79 net79 clock_out[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2842__D u1.col_sel\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1908__A1 _0360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3077__CLK clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1480_ u1.ordering_timer\[15\] _1097_ u1.ordering_timer\[11\] _1104_ _1105_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3150_ net47 net72 spi_data_crossing\[16\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3081_ _0007_ clknet_leaf_9_clock u0.run_state\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2078__S _0470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2101_ _0457_ _0490_ _0492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3261__I clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2032_ _0443_ _0076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2914__CLK clknet_leaf_7_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2934_ _0076_ clknet_leaf_28_clock u1.ccr1\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2865_ reset_n clknet_leaf_37_clock reset_n_sync\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1816_ net37 _1144_ _0293_ _0001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2796_ u1.ccr0\[3\] _0363_ _1013_ _1020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1747_ _1207_ _1364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1678_ u1.timer\[10\] _1295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3279_ net110 net126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2937__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1841__A3 _1155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2650_ _1266_ _0908_ _0910_ _0917_ _0918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_12_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1601_ _1213_ u1.timer\[3\] _1219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3256__I clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2581_ _0863_ _0205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2160__I _0528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2554__A1 _0447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1532_ u0.run_state\[0\] _1154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2554__B2 spi_data_crossing\[16\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1463_ u1.ordering_timer\[25\] _1088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3202_ _0272_ clknet_leaf_7_clock u1.ccr0\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input1_I io_control_trigger_in vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3133_ spi_data_crossing\[7\].A clknet_leaf_2_clock spi_data_crossing\[7\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3064_ _0206_ clknet_leaf_12_clock u0.cmd\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2015_ u1.ccr1\[21\] _0367_ _0427_ _0434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1832__A3 _0296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3242__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2917_ _0059_ clknet_leaf_4_clock u1.ccr1\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2848_ u0.cmd\[4\] clknet_leaf_23_clock net105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2779_ net5 _1008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input57_I spi_data[25] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_9_clock_I clknet_2_1__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2784__A1 _0447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1587__A2 _1204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2536__A1 _0379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3115__CLK clknet_leaf_29_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2075__I0 _0474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2702_ _1295_ _0956_ _0960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2633_ latch_data_sync\[0\] latch_data latch_data_sync\[1\] _1042_ _0904_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and4_1
Xoutput214 net214 row_select_right[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput203 net203 row_col_select[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2564_ u0.cmd\[20\] _0852_ _0853_ spi_data_crossing\[20\].data_sync _0854_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1515_ u1.ordering_timer\[1\] _1134_ _1140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2495_ _1082_ _0801_ _0805_ _0806_ _0725_ _0807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_1446_ u1.ordering_timer\[28\] _1071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1502__A2 _1126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3116_ _0250_ clknet_leaf_29_clock u1.timer\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3047_ _0189_ clknet_leaf_3_clock u0.cmd\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1813__I0 net18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2518__B2 spi_data_crossing\[3\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2518__A1 _0462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output163_I net163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3138__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2850__D u0.cmd\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2509__A1 _1042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2280_ u1.ordering_timer\[3\] _0612_ _0619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_42_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2460__A3 _0776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1995_ _1253_ _0416_ _0420_ _0062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2748__A1 _0983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2613__I _0890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2616_ _0891_ _0892_ _0893_ _0210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_47_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2547_ _0842_ _0192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1723__A2 _1337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2478_ _1093_ _0790_ _0791_ _0792_ _0793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1429_ u1.ordering_complete\[23\] _1054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output88_I net88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2211__I0 _0365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2845__D u0.cmd\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1780_ _1395_ _1396_ _1359_ _1397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2202__I0 _0513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2401_ _1068_ _0721_ _0724_ _0725_ _0726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2332_ _0648_ u1.ordering_timer\[9\] _0654_ _0649_ _0665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_27_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2263_ _0603_ _0604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2194_ _0472_ u1.inverter_select\[7\] _0545_ _0549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1469__B2 u1.ordering_complete\[26\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1469__A1 _1093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_36_clock_I clknet_2_0__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2418__B1 _0734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1978_ _0372_ _0407_ _0411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1944__A2 _0378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2970__CLK clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2657__B1 _1235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2672__A3 _1204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1880__A1 _0330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_15_clock clknet_2_1__leaf_clock clknet_leaf_15_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1935__A2 _0378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2360__A2 _0682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2950_ _0092_ clknet_leaf_4_clock u1.ordering_complete\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3259__I clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2881_ _0015_ clknet_leaf_11_clock u0.mem_write_n\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1901_ u0.cmd\[1\] _0356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1832_ _0299_ _1160_ _0296_ _0302_ _0015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2843__CLK clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1763_ _1289_ _1290_ _1379_ _1380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1694_ _1262_ _1311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2993__CLK clknet_leaf_22_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3295_ net148 net147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2315_ _1124_ _0649_ _0650_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2246_ _1057_ _0584_ _0586_ _0587_ _1055_ _0588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__2338__I _0610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2177_ u0.cmd\[19\] _0350_ _0448_ _0539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_41_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1614__A1 _1227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2590__A2 _0864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1417__I _1041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2342__A2 _0655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2866__CLK clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1908__A2 _0361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2333__A2 _0665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3080_ _0005_ clknet_leaf_12_clock u0.run_state\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2100_ _1060_ _0489_ _0491_ _0096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2031_ u1.ccr1\[28\] _0442_ _0438_ _0443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_0 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2933_ _0075_ clknet_leaf_25_clock u1.ccr1\[27\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2864_ control_trigger_sync\[0\] clknet_leaf_15_clock control_trigger_sync\[1\] vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2795_ _1019_ _0263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1815_ net19 net37 _0293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1746_ _1209_ _1363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3021__CLK clknet_leaf_35_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1677_ _1269_ u1.ccr0\[11\] u1.ccr0\[10\] _1268_ _1294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__3171__CLK clknet_leaf_10_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1681__B _1297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3278_ net109 net125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2068__I _0451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2229_ _1096_ _0571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1835__A1 _0298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2889__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_5_clock_I clknet_2_0__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2012__A1 _0429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2531__I _0820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2687__B _1280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1811__S net35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2853__D u0.cmd\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3044__CLK clknet_leaf_7_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1600_ u1.ccr1\[1\] _1209_ _1218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2580_ _1160_ _0858_ _0859_ spi_data_crossing\[27\].data_sync _0863_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3194__CLK clknet_leaf_16_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1531_ u0.cmd\[29\] _1153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2597__B _1212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1462_ u1.ordering_timer\[26\] _1087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__3272__I net103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3201_ _0271_ clknet_leaf_3_clock u1.ccr0\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3132_ net69 net72 spi_data_crossing\[7\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3063_ _0205_ clknet_leaf_11_clock u0.cmd\[27\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1817__A1 u0.cmd\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2014_ _0433_ _0068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1520__I _1144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2490__A1 u1.ordering_complete\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2916_ _0058_ clknet_leaf_3_clock u1.ccr1\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2847_ u0.cmd\[3\] clknet_leaf_19_clock net104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2778_ _1007_ net24 _0258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1729_ _1177_ _1343_ _1344_ _1345_ _1346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1505__B1 _1122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3067__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2481__A1 _1093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2904__CLK clknet_leaf_28_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2848__D u0.cmd\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2472__A1 _0711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2224__A1 _1070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2075__I1 _1112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2701_ _1295_ _0956_ _0959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2632_ _0891_ _0903_ _0216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput204 net204 row_select_left[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput215 net215 row_select_right[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2563_ _0846_ _0853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1514_ _1138_ _1139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2494_ u1.ordering_timer\[28\] _0791_ _0806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1445_ _1057_ _1063_ _1066_ _1069_ _1070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3115_ _0249_ clknet_leaf_29_clock u1.timer\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3046_ _0188_ clknet_leaf_3_clock u0.cmd\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2463__A1 _0774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2927__CLK clknet_leaf_23_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1569__A3 _1182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1813__I1 net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2454__A1 _0735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2509__A2 u0.latch_cmd vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3232__CLK clknet_leaf_22_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2367__S _0607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1994_ _0387_ _0394_ _0420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1420__A2 _1044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_32_clock_I clknet_2_2__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2615_ u1.row_sel\[0\] _0875_ _0893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2546_ _0387_ _0838_ _0839_ spi_data_crossing\[14\].data_sync _0842_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1723__A3 _1338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2477_ _0725_ _0792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1428_ _1047_ u1.ordering_complete\[22\] _1049_ u1.ordering_complete\[21\] _1053_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_28_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3029_ _0171_ clknet_leaf_30_clock u1.ordering_timer\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2436__A1 _1047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3105__CLK clknet_leaf_26_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2675__A1 _1214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2861__D latch_data vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ _0596_ _0725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2331_ _1109_ _0663_ _0664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2262_ _0602_ _0603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3280__I net96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2193_ _0548_ _0132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1469__A2 u1.ordering_complete\[27\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3128__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1977_ _1200_ _0409_ _0410_ _0054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2529_ _0831_ _0185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input32_I la_oenb[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2657__B2 _0923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2409__A1 _0329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2196__I0 _0474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1699__A2 _1308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2856__D u0.cmd\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2120__I0 _0476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2880_ _0014_ clknet_leaf_11_clock u0.mem_write_n\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1900_ _0355_ _0032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2820__A1 u0.cmd\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1831_ _0296_ _0302_ _0303_ _0014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_42_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2584__B1 _0865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1762_ _1284_ _1288_ _1291_ _1379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3275__I net106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1693_ u1.ccr0\[12\] _1310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2336__B1 _0662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3294_ net146 net145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2314_ u1.ordering_timer\[6\] u1.ordering_timer\[5\] _0623_ _0627_ _0649_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2245_ _1051_ _1053_ _1048_ _0587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2176_ _0310_ _0530_ _0538_ _0125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2111__I0 _0466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_1_clock_I clknet_2_0__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2566__B1 _0853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2169__I0 _0462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2030_ u0.cmd\[12\] _0442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_2932_ _0074_ clknet_leaf_25_clock u1.ccr1\[26\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2863_ control_trigger clknet_leaf_15_clock control_trigger_sync\[0\] vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2794_ u1.ccr0\[2\] _0360_ _1017_ _1019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1814_ _0292_ _0000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2960__CLK clknet_leaf_33_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1745_ _1347_ _1356_ _1361_ _1362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_11_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1676_ u1.timer\[9\] _1293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3277_ net108 net124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2228_ _1132_ _0568_ _0569_ _1129_ _0570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1835__A2 _0305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2159_ _0447_ _0348_ _0450_ _0528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_26_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_14_clock clknet_2_1__leaf_clock clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_26_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_29_clock clknet_2_2__leaf_clock clknet_leaf_29_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_6_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output186_I net186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2012__A2 _0430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2833__CLK clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2983__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1530_ _1043_ _1152_ _0008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1461_ u1.ordering_complete\[24\] _1086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3200_ _0270_ clknet_leaf_27_clock u1.ccr0\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3131_ spi_data_crossing\[6\].A clknet_leaf_0_clock spi_data_crossing\[6\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3062_ _0204_ clknet_leaf_11_clock u0.cmd\[26\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2013_ u1.ccr1\[20\] _0365_ _0427_ _0433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2490__A2 _0720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2915_ _0057_ clknet_leaf_3_clock u1.ccr1\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2846_ u0.cmd\[2\] clknet_leaf_17_clock net103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2777_ net6 _1007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1753__A1 _1204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1728_ u1.timer\[26\] _1345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1659_ _1251_ _1266_ _1276_ _1277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2856__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1505__A1 _1128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1808__A2 _1403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_27_clock_I clknet_2_2__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output101_I net101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2481__A2 _0710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1867__B _0329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1992__A1 u0.cmd\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3011__CLK clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3161__CLK clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2224__A2 _1095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2700_ _0945_ _0958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1983__A1 u0.cmd\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2631_ u1.row_sel\[5\] _0900_ u1.row_sel\[6\] _0903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput205 net205 row_select_left[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2562_ _0844_ _0852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2879__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3283__I net99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2401__B _0724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1513_ u1.ordering_timer\[0\] _1138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2493_ _1082_ u1.ordering_timer\[29\] _0805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1444_ u1.ordering_timer\[18\] _1067_ _1068_ _1061_ _1069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_3114_ _0248_ clknet_leaf_29_clock u1.timer\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1531__I u0.cmd\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3045_ _0187_ clknet_leaf_3_clock u0.cmd\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2463__A2 _0779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2362__I _0634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1423__B1 _1047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1974__A1 _1196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2829_ _1038_ _0278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input62_I spi_data[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3034__CLK clknet_leaf_33_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2151__A1 _0404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3184__CLK clknet_leaf_36_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2859__D u0.cmd\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1717__B2 _1237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1717__A1 _1236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2693__A2 _0951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3278__I net109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1993_ _1263_ _0416_ _0419_ _0061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2614_ u1.row_sel\[0\] _0875_ _0892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3057__CLK clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2545_ _0841_ _0191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2476_ u1.ordering_timer\[27\] _0783_ _1085_ _0784_ _0791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1427_ _1048_ _1051_ _1052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2133__A1 u0.cmd\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2357__I _0629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3028_ _0170_ clknet_leaf_31_clock u1.ordering_timer\[24\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2436__A2 _0750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1947__A1 _1353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2124__A1 _0504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2330_ _0654_ _0656_ _0663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2261_ _0565_ _0600_ _0602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2917__CLK clknet_leaf_4_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2192_ _0469_ u1.inverter_select\[6\] _0545_ _0548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2418__A2 _0719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1976_ _0369_ _0407_ _0410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2528_ _0472_ _0826_ _0827_ spi_data_crossing\[7\].data_sync _0831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2459_ _0676_ _1116_ _0775_ _0692_ _0776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__2106__A1 _0402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input25_I la_oenb[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2815__I u1.ccr0\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3222__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2196__I1 u1.inverter_select\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2198__S _0539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1699__A3 _1309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3033__D _0175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1769__C _1385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2120__I1 u1.ordering_complete\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2820__A2 _1029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1830_ u0.cmd\[26\] _1149_ _0303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1761_ _1292_ _1369_ _1378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1692_ _1293_ u1.ccr0\[9\] u1.ccr0\[8\] _1267_ _1309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_48_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2313_ u1.ordering_timer\[7\] _0648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1804__I u1.timer\[22\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3293_ net144 net143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2244_ _1066_ _0585_ _0586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2175_ _0468_ _0531_ _0538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3245__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2111__I1 u1.ordering_complete\[21\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1959_ _0393_ _0397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2370__I u1.ordering_timer\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2802__A2 _1014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2566__A1 u0.cmd\[21\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2566__B2 spi_data_crossing\[21\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2318__A1 _0648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3118__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2867__D _0024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2931_ _0073_ clknet_leaf_27_clock u1.ccr1\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2862_ latch_data_sync\[0\] clknet_leaf_7_clock latch_data_sync\[1\] vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2793_ _1018_ _0262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1813_ net18 net1 net36 _0292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1744_ _1359_ _1360_ _1361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1675_ _1285_ _1288_ _1291_ _1292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2309__A1 u1.ordering_complete\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3276_ net107 net123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2227_ _1123_ _1131_ _1126_ _0569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2158_ _0526_ _0522_ _0527_ _0118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2365__I _0693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2089_ u0.cmd\[14\] _0478_ _0483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_23_clock_I clknet_2_3__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2548__B2 spi_data_crossing\[15\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2548__A1 _0389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1523__A2 control_trigger vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2720__A1 _0283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2087__I0 _0385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1460_ u1.ordering_timer\[24\] _1085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3090__CLK clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3130_ net68 net72 spi_data_crossing\[6\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2711__A1 _0935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3061_ _0203_ clknet_leaf_11_clock u0.cmd\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1817__A3 _1155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2012_ _0429_ _0430_ _0432_ _0067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2078__I0 _0476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2914_ _0056_ clknet_leaf_7_clock u1.ccr1\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2845_ u0.cmd\[1\] clknet_leaf_18_clock net102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1450__B2 u1.ordering_complete\[27\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2776_ _1006_ net25 _0257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1727_ u1.ccr0\[26\] _1344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1753__A2 u1.ccr0\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1658_ u1.ccr1\[8\] _1267_ _1274_ _1275_ _1276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1589_ _1206_ _1207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1505__A2 u1.ordering_complete\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3259_ clknet_leaf_12_clock net78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2095__I _0486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2069__I0 _0469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1992__A2 _0413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2792__I1 _0356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2950__CLK clknet_leaf_4_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2630_ _0891_ _0902_ _0215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1983__A2 _0413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput206 net206 row_select_left[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2561_ _0851_ _0197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_13_clock clknet_2_1__leaf_clock clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2492_ u1.ordering_complete\[30\] _0792_ _0804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1512_ _1128_ u1.ordering_complete\[3\] _1136_ u1.ordering_complete\[2\] _1137_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_1443_ u1.ordering_timer\[17\] _1068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2401__C _0725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3216__D u1.inverter_select\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3113_ _0247_ clknet_leaf_24_clock u1.timer\[27\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1812__I _0291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_28_clock clknet_2_2__leaf_clock clknet_leaf_28_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3044_ _0186_ clknet_leaf_7_clock u0.cmd\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1671__A1 _1283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1974__A2 _0398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1423__B2 u1.ordering_complete\[22\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2828_ net13 net31 _1038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2759_ _0996_ _0995_ _0997_ _0934_ _0249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_30_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input55_I spi_data[23] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2973__CLK clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3036__D _0178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2875__D u0.latch_cmd vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2846__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1992_ u0.cmd\[13\] _0413_ _0419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2613_ _0890_ _0891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3294__I net146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2996__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2544_ _0385_ _0838_ _0839_ spi_data_crossing\[13\].data_sync _0841_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2475_ _0783_ _0774_ _0779_ _0790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1426_ _1049_ u1.ordering_complete\[21\] _1050_ u1.ordering_complete\[20\] _1051_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_25_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2133__A2 _0507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3027_ _0169_ clknet_leaf_32_clock u1.ordering_timer\[23\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1947__A2 _0361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3001__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2372__A2 _0687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3151__CLK clknet_leaf_7_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2124__A2 _0500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1883__A1 _0330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2869__CLK clknet_leaf_18_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1938__A2 _0378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2260_ _0600_ _0601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2191_ _0547_ _0131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1874__A1 _0331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1975_ _0397_ _0409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3024__CLK clknet_leaf_32_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2051__A1 _0457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3174__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2527_ _0830_ _0184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2458_ _0648_ u1.ordering_timer\[9\] _0654_ _0649_ _0775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_29_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2106__A2 _0493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2389_ u1.ordering_complete\[16\] _0714_ _0715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input18_I la_data_in[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2290__A1 _1122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1447__I u1.ordering_timer\[27\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_2_2__f_clock clknet_0_clock clknet_2_2__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1910__I u0.cmd\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_18_clock_I clknet_2_3__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2227__B _1126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3047__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2281__A1 u1.ordering_complete\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1760_ _1370_ _1376_ _1368_ _1377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2584__A2 _0864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3197__CLK clknet_leaf_15_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1691_ _1306_ _1307_ _1308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2336__A2 _0655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2312_ _0647_ _0152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3292_ net142 net141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2243_ _1062_ _1069_ _0585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2174_ _0537_ _0124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2272__A1 _1138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1958_ _0396_ _0049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1889_ u0.cmd\[0\] _0345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2327__A2 _0655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1838__A1 _0299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2907__CLK clknet_leaf_15_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2566__A2 _0852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2810__I0 u1.ccr0\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2002__S _0423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1905__I _0358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2883__D _0017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1640__I u1.timer\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2930_ _0072_ clknet_leaf_25_clock u1.ccr1\[24\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2861_ latch_data clknet_leaf_2_clock latch_data_sync\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2792_ u1.ccr0\[1\] _0356_ _1017_ _1018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1812_ _0291_ _0002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1743_ _1167_ u1.ccr0\[30\] u1.ccr0\[29\] _1168_ _1360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1674_ _1289_ _1290_ _1281_ _1280_ _1291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1765__B1 _1299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2309__A2 _0630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3275_ net106 net122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3212__CLK clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2226_ _1141_ _0567_ _1137_ _0568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2157_ _0468_ _0515_ _0527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2493__A1 _1082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1550__I u1.timer\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2088_ _0482_ _0093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2484__A1 _0597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2087__I1 u1.ordering_complete\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2878__D _0012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3235__CLK clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3060_ _0202_ clknet_leaf_11_clock u0.cmd\[24\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2011_ _0402_ _0431_ _0432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2078__I1 _1110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3297__I net163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2913_ _0055_ clknet_leaf_7_clock u1.ccr1\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2844_ u0.cmd\[0\] clknet_leaf_17_clock net95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1450__A2 u1.ordering_complete\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2775_ net7 _1006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1738__B1 u1.ccr0\[24\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1726_ u1.ccr0\[27\] _1343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1545__I u1.timer\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1657_ _1247_ _1248_ _1275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2002__I1 _0356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1588_ u1.timer\[0\] _1206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3258_ clknet_leaf_12_clock net77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2376__I _1096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2209_ _0557_ _0139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3189_ _0259_ clknet_leaf_37_clock net153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3108__CLK clknet_leaf_24_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2069__I1 u1.ordering_complete\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1729__B1 _1344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_9_clock clknet_2_1__leaf_clock clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1680__A2 u1.ccr0\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2235__B _0573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput207 net207 row_select_left[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2560_ u0.cmd\[19\] _0845_ _0847_ spi_data_crossing\[19\].data_sync _0851_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2491_ _1076_ _0709_ _0803_ _0565_ _0175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1511_ u1.ordering_timer\[2\] _1136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1442_ u1.ordering_complete\[18\] _1067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3112_ _0246_ clknet_leaf_24_clock u1.timer\[26\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3232__D u1.row_col_select\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3043_ _0185_ clknet_leaf_2_clock u0.cmd\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2827_ _1037_ _0277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2758_ _0996_ _0995_ _0997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1709_ _1324_ _1325_ _1326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2689_ u1.timer\[7\] u1.timer\[4\] _0941_ _0947_ _0950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA_input48_I spi_data[17] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2687__A1 _1283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2439__A1 _0735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3080__CLK clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1913__I u0.cmd\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1991_ _1261_ _0416_ _0418_ _0060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2612_ _0875_ _0889_ _0890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_16_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2543_ _0840_ _0190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3227__D u1.row_col_select\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2474_ _0789_ _0172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2669__A1 _1364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1425_ u1.ordering_timer\[20\] _1050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3026_ _0168_ clknet_leaf_31_clock u1.ordering_timer\[22\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2940__CLK clknet_leaf_4_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3137__D spi_data_crossing\[9\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1580__A1 _1196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1580__B2 u1.timer\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2829__I _1038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_12_clock clknet_2_1__leaf_clock clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_14_clock_I clknet_2_1__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_27_clock clknet_2_2__leaf_clock clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_6_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2190_ _0367_ u1.inverter_select\[5\] _0545_ _0547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2474__I _0789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1974_ _1196_ _0398_ _0408_ _0053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2963__CLK clknet_leaf_30_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2051__A2 _0455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2526_ _0469_ _0826_ _0827_ spi_data_crossing\[6\].data_sync _0830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2457_ u1.ordering_timer\[25\] _0774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2388_ _0606_ _0714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_29_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3009_ _0151_ clknet_leaf_0_clock u1.ordering_timer\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2384__I _0709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2814__A1 _1296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2290__A2 _0627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2042__A2 u0.cmd\[21\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1728__I u1.timer\[26\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2836__CLK clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2986__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2281__A2 _0597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1638__I u1.timer\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1792__A1 _1406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1690_ _1256_ u1.ccr0\[15\] u1.ccr0\[14\] _1257_ _1307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1544__A1 _1043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2311_ u1.ordering_timer\[6\] _0626_ _0635_ _0646_ _0647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3291_ net140 net139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2242_ _0583_ _1058_ _0584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2173_ _0466_ u1.col_limit\[5\] _0529_ _0537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1480__B1 u1.ordering_timer\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3141__CLK clknet_leaf_2_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1957_ u1.ccr1\[1\] _0356_ _0394_ _0396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1548__I _1165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1888_ _0331_ _0344_ _0031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1783__A1 _1362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2859__CLK clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2509_ _1042_ u0.latch_cmd _0819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input30_I la_oenb[17] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1838__A2 _1160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2810__I1 _0376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3014__CLK clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3164__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2860_ u1.output_active clknet_leaf_7_clock net192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1811_ net17 net2 net35 _0291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2791_ _1012_ _1017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1765__A1 _1294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1742_ u1.timer\[29\] _1357_ _1358_ u1.timer\[28\] _1359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1673_ u1.ccr0\[7\] _1290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1765__B2 _1309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3235__D u0.cmd\[17\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3274_ net105 net121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2225_ _1135_ _1140_ _0567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2156_ u1.row_limit\[6\] _0526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2493__A2 u1.ordering_timer\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2087_ _0385_ u1.ordering_complete\[13\] _0452_ _0482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2989_ _0131_ clknet_leaf_22_clock u1.inverter_select\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1756__A1 _1362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3037__CLK clknet_leaf_15_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3187__CLK clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1692__B1 u1.ccr0\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2236__A2 _0577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1444__B1 _1068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1916__I u0.cmd\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2013__S _0427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2010_ _0422_ _0431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2475__A2 _0774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2227__A2 _1131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2912_ _0054_ clknet_leaf_7_clock u1.ccr1\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2843_ u1.col_sel\[5\] clknet_leaf_19_clock net88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2774_ _1005_ net26 _0256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1725_ _1323_ _1326_ _1341_ _1342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1738__A1 _1171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1656_ u1.ccr1\[10\] _1268_ _1270_ _1273_ _1274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1587_ u1.ccr1\[2\] _1204_ _1205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2163__A1 _0454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3257_ clknet_leaf_12_clock net76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2208_ _0363_ u1.row_col_select\[3\] _0553_ _0557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3188_ _0258_ clknet_leaf_37_clock net155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2139_ _0514_ _0515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1977__A1 _1200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1729__B2 _1345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2154__A1 _0406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1471__I u1.ordering_timer\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3202__CLK clknet_leaf_7_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput208 net208 row_select_left[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_12_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2490_ u1.ordering_complete\[29\] _0720_ _0709_ _0802_ _0803_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1510_ u1.ordering_timer\[0\] _1133_ u1.ordering_timer\[1\] _1134_ _1135_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_4_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1441_ _1064_ u1.ordering_complete\[19\] _1065_ u1.ordering_complete\[18\] _1066_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_3111_ _0245_ clknet_leaf_29_clock u1.timer\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2477__I _0725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2696__A2 _1267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3042_ _0184_ clknet_leaf_7_clock u0.cmd\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2448__A2 _0720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2826_ net4 net22 _1037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_20_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2757_ u1.timer\[29\] _0996_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1708_ _1318_ _1319_ _1325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2688_ _0946_ _0948_ _0949_ _0226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1639_ u1.timer\[14\] _1257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2136__A1 _1073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2687__A2 _0942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3309_ net206 net212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3225__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2127__A1 u0.cmd\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2678__A2 _0941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2297__I _0602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_10_clock_I clknet_2_1__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1990_ u0.cmd\[12\] _0413_ _0418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2611_ _0886_ _0887_ _0888_ _0329_ _0889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_6_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2542_ _0442_ _0838_ _0839_ spi_data_crossing\[12\].data_sync _0840_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2473_ _0783_ _0716_ _0762_ _0788_ _0789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2892__CLK clknet_leaf_26_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1424_ u1.ordering_timer\[21\] _1049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3248__CLK clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3025_ _0167_ clknet_leaf_32_clock u1.ordering_timer\[21\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_8_clock clknet_2_1__leaf_clock clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_20_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2809_ _1027_ _0269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input60_I spi_data[28] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1955__I1 _0345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2111__S _0496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2021__S _0427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1859__B1 u1.col_sel\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2823__A2 _1015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1973_ _0406_ _0407_ _0408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3238__D u0.cmd\[20\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2525_ _0829_ _0183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2456_ _0773_ _0170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3070__CLK clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2387_ _1059_ _0712_ _0713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3008_ _0150_ clknet_leaf_1_clock u1.ordering_timer\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2814__A2 _1025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2578__A1 _0299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2578__B2 spi_data_crossing\[26\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2042__A3 u0.cmd\[20\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1919__I u0.cmd\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3093__CLK clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3290_ net157 net156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2310_ _0643_ _0644_ _0645_ _0646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2241_ u1.ordering_timer\[19\] _0583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2172_ _0536_ _0123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2930__CLK clknet_leaf_25_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1480__B2 _1104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1480__A1 u1.ordering_timer\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1956_ _0395_ _0048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1887_ u1.col_sel\[6\] _0343_ _0344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2508_ _0817_ _0818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2732__A1 _0937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_11_clock clknet_2_1__leaf_clock clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2439_ _0735_ _0756_ _0758_ _0759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input23_I la_oenb[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_26_clock clknet_2_3__leaf_clock clknet_leaf_26_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_29_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2395__I _0610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2799__A1 _0404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output91_I net91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2723__A1 _0282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2953__CLK clknet_leaf_35_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1810_ _0290_ _0003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2790_ _1010_ _1014_ _1016_ _0261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1741_ u1.ccr0\[28\] _1358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1765__A2 _1297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1672_ u1.timer\[7\] _1289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2714__A1 _0958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3273_ net104 net120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2224_ _1070_ _1095_ _0566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2155_ _0524_ _0522_ _0525_ _0117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2086_ _0481_ _0092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1559__I u1.timer\[27\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2988_ _0130_ clknet_leaf_22_clock u1.inverter_select\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1939_ _0353_ _0383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2611__C _0329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2976__CLK clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2705__A1 _1272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1692__B2 _1267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1444__B2 _1061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1995__A2 _0416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1932__I _0358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3131__CLK clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2475__A3 _0779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2849__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2911_ _0053_ clknet_leaf_7_clock u1.ccr1\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2842_ u1.col_sel\[4\] clknet_leaf_19_clock net87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2773_ net8 _1005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2999__CLK clknet_leaf_22_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1724_ _1333_ _1334_ _1335_ _1340_ _1341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__1738__A2 u1.ccr0\[31\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1655_ _1271_ _1272_ u1.ccr1\[10\] _1268_ _1273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1586_ _1203_ _1204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3256_ clknet_leaf_12_clock net75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2207_ _0556_ _0138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3187_ _0257_ clknet_leaf_37_clock net157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2138_ _0346_ _0348_ _0450_ _0514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__1674__B2 _1280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2069_ _0469_ u1.ordering_complete\[6\] _0470_ _0471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1426__B2 u1.ordering_complete\[20\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3004__CLK clknet_leaf_34_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3154__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2217__I0 _0472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2024__S _0438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2393__A2 _0710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput209 net209 row_select_left[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_4_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1440_ u1.ordering_timer\[18\] _1065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1662__I _1279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3110_ _0244_ clknet_leaf_24_clock u1.timer\[24\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3041_ _0183_ clknet_leaf_7_clock u0.cmd\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1656__A1 u1.ccr1\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2605__B1 u1.row_limit\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3027__CLK clknet_leaf_32_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2081__A1 u0.cmd\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2208__I0 _0363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2825_ _1304_ _1015_ _1036_ _0276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3177__CLK clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2756_ _0982_ _0994_ _0995_ _0248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1707_ _1321_ _1320_ _1324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2687_ _1283_ _0942_ _1280_ _0949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1592__B1 u1.ccr1\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1638_ u1.timer\[15\] _1256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2136__A2 _0490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1569_ _1170_ _1175_ _1182_ _1186_ _1187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3308_ net205 net211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1505__C _1129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3239_ u0.cmd\[21\] clknet_leaf_9_clock net167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1647__A1 _1261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2109__S _0496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1583__B1 _1200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2127__A2 _0507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2610_ u1.row_sel\[6\] _0526_ _0888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2541_ _0820_ _0839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2472_ _0711_ _0786_ _0787_ _0788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1423_ _1046_ u1.ordering_complete\[23\] _1047_ u1.ordering_complete\[22\] _1048_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1877__A1 _0330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3024_ _0166_ clknet_leaf_32_clock u1.ordering_timer\[20\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2808_ u1.ccr0\[8\] _0374_ _1013_ _1027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2739_ _0286_ _0981_ _0985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_3_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input53_I spi_data[21] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2348__A2 _0658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1556__B1 u1.ccr1\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1859__B2 _0318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2771__I net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1972_ _0393_ _0407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2339__A2 _0665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2524_ _0466_ _0826_ _0827_ spi_data_crossing\[5\].data_sync _0829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3215__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2455_ _0769_ _0755_ _0762_ _0772_ _0773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2386_ _0703_ _0698_ _0694_ _0712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_29_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3007_ _0149_ clknet_leaf_4_clock u1.ordering_timer\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2882__CLK clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3238__CLK clknet_leaf_10_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2240_ _1202_ _1277_ _0579_ _0581_ _0582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_26_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2171_ _0464_ u1.col_limit\[4\] _0529_ _0536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1670__I u1.timer\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_7_clock clknet_2_1__leaf_clock clknet_leaf_7_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_24_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2257__A1 _0565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1955_ u1.ccr1\[0\] _0345_ _0394_ _0395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1886_ u1.col_sel\[5\] _0340_ _0343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2507_ _0816_ _0817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2438_ u1.ordering_complete\[22\] _0757_ _0758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2369_ _0697_ _0159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1838__A4 _0305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input16_I la_data_in[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2248__A1 _1084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2799__A2 _1021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3300__I net166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2487__A1 u1.ordering_timer\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3060__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1740_ u1.ccr0\[29\] _1357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1671_ _1283_ _1282_ _1286_ _1287_ _1288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2714__A2 _0966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3272_ net103 net119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I la_data_in[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2478__A1 _1093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2223_ _1402_ _0565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_23_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2154_ _0406_ _0515_ _0525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2085_ _0442_ u1.ordering_complete\[12\] _0452_ _0481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2650__A1 _1266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2987_ _0129_ clknet_leaf_19_clock u1.inverter_select\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1938_ _1343_ _0378_ _0382_ _0043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2402__A1 _1061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1869_ _1212_ _0309_ _0332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1575__I u1.timer\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2469__A1 _0769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1692__A2 u1.ccr0\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3083__CLK clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1485__I u1.ordering_complete\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2920__CLK clknet_leaf_33_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2632__A1 _0891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2910_ _0052_ clknet_leaf_6_clock u1.ccr1\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_10_clock clknet_2_1__leaf_clock clknet_leaf_10_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_32_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2841_ u1.col_sel\[3\] clknet_leaf_19_clock net86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2772_ _1004_ net27 _0255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1723_ _1336_ _1337_ _1338_ _1339_ _1340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xclkbuf_leaf_25_clock clknet_2_3__leaf_clock clknet_leaf_25_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1654_ u1.timer\[11\] _1272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1585_ u1.timer\[2\] _1203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2699__A1 _0946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3255_ clknet_leaf_12_clock net74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2206_ _0360_ u1.row_col_select\[2\] _0553_ _0556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2171__I0 _0464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3186_ _0256_ clknet_leaf_36_clock net140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2137_ _0454_ _0513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1674__A2 _1290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2068_ _0451_ _0470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_41_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1426__A2 u1.ordering_complete\[21\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2943__CLK clknet_leaf_1_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1985__I0 u1.ccr1\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2614__A1 u1.row_sel\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2090__A2 _0455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3040_ _0182_ clknet_leaf_8_clock u0.cmd\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1656__A2 _1268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2605__A1 u1.row_limit\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2966__CLK clknet_leaf_28_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2081__A2 _0478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2215__S _0558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2208__I1 u1.row_col_select\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2824_ u0.cmd\[15\] _1017_ _1036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2755_ _1413_ _0993_ _0995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1706_ _1318_ _1319_ _1320_ _1322_ _1323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_2686_ _0942_ _0947_ _0948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1853__I u1.col_sel\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1637_ _1252_ u1.timer\[15\] _1253_ _1254_ _1255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3307_ net204 net210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1568_ _1183_ _1184_ _1185_ _1186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1499_ u1.ordering_timer\[7\] _1124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3238_ u0.cmd\[20\] clknet_leaf_10_clock net166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3169_ spi_data_crossing\[25\].A clknet_leaf_10_clock spi_data_crossing\[25\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2684__I _0945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3121__CLK clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1583__A1 _1199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2839__CLK clknet_leaf_18_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2989__CLK clknet_leaf_22_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2035__S _0438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2540_ _0817_ _0838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1574__A1 u1.ccr1\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1673__I u1.ccr0\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2769__I net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2471_ u1.ordering_complete\[26\] _0757_ _0787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1422_ u1.ordering_timer\[22\] _1047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_37_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3023_ _0165_ clknet_leaf_36_clock u1.ordering_timer\[19\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2826__A1 net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2009__I _0426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3144__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2807_ _1290_ _1025_ _1026_ _0268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2738_ _0286_ _0981_ _0984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1565__A1 u1.ccr1\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2669_ _1364_ _1208_ _0936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_8_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input46_I spi_data[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3303__I net169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2293__A2 _0630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1556__B2 _1173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1556__A1 u1.ccr1\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1859__A2 _0321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3017__CLK clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3167__CLK clknet_leaf_10_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1492__B1 _1109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1971_ u0.cmd\[5\] _0406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1795__A1 _1394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2499__I u1.ordering_timer\[31\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2523_ _0828_ _0182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2454_ _0735_ _0770_ _0771_ _0772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2385_ _0606_ _0711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput1 io_control_trigger_in net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3006_ _0148_ clknet_leaf_4_clock u1.ordering_timer\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2027__A2 _0430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1786__A1 _1402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1474__B1 u1.ordering_timer\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2018__A2 _0430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2821__B _1034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1951__I u0.cmd\[17\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2170_ _0535_ _0122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1954_ _0393_ _0394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_21_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1885_ _0331_ _0342_ _0030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2506_ _0815_ u0.latch_cmd _0816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2437_ _0629_ _0757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1940__A1 u0.cmd\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2368_ u1.ordering_timer\[13\] _0682_ _0691_ _0696_ _0697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2299_ u1.ordering_timer\[5\] _0623_ _0627_ _0636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_38_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1759__A1 _1363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2420__A2 _0737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3175__D spi_data_crossing\[28\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2723__A3 _0970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput190 net190 mem_write_n[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2487__A2 _0791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1695__B1 _1310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3205__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1670_ u1.timer\[4\] _1287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3085__D _0219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2175__A1 _0468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2777__I net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3271_ net102 net118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2222_ _0564_ _0145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2153_ u1.row_limit\[5\] _0524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2084_ _1104_ _0453_ _0480_ _0091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_19_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1438__B1 _1059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2986_ _0128_ clknet_leaf_20_clock u1.inverter_select\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1937_ _0381_ _0370_ _0382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2402__A2 _0720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1868_ _0330_ _0331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput70 spi_data[8] net70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2166__A1 _0318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1799_ _1318_ _0281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2872__CLK clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2469__A2 _0784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1677__B1 u1.ccr0\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3228__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2641__A2 _1303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_6_clock clknet_2_1__leaf_clock clknet_leaf_6_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_5_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2157__A1 _0468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2840_ u1.col_sel\[2\] clknet_leaf_18_clock net85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2771_ net9 _1004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1722_ _1237_ u1.ccr0\[16\] _1339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1653_ u1.ccr1\[11\] _1271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2895__CLK clknet_leaf_23_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1584_ _1192_ _1195_ _1198_ _1201_ _1202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3254_ clknet_leaf_12_clock net73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2205_ _0555_ _0137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2171__I1 u1.col_limit\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3185_ _0255_ clknet_leaf_36_clock net142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2136_ _1073_ _0490_ _0512_ _0111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2067_ _0468_ _0469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2969_ _0111_ clknet_leaf_28_clock u1.ordering_complete\[31\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2387__A1 _1059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1985__I1 _0379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3306__I net192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2210__I _0552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2311__A1 u1.ordering_timer\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3050__CLK clknet_leaf_4_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2366__B _0694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2614__A2 _0875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2823_ _1305_ _1015_ _1035_ _0275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2754_ _1413_ _0993_ _0994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1705_ _1321_ _1322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2685_ u1.timer\[6\] u1.timer\[5\] _0947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1636_ u1.timer\[14\] _1254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3073__CLK clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1567_ u1.ccr1\[31\] _1171_ _1185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3306_ net192 net193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2030__I u0.cmd\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1498_ _1121_ u1.ordering_complete\[5\] _1122_ u1.ordering_complete\[4\] _1123_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3237_ u0.cmd\[19\] clknet_leaf_9_clock net165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3168_ net57 net72 spi_data_crossing\[25\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2119_ _0502_ _0104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2910__CLK clknet_leaf_6_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3099_ _0233_ clknet_leaf_27_clock u1.timer\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1583__A2 u1.timer\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2780__A1 _1008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3183__D _0253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2532__A1 _0474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_24_clock clknet_2_3__leaf_clock clknet_leaf_24_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_18_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2115__I _0488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1954__I _0393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3096__CLK clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2470_ _1087_ _0785_ _0786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1421_ u1.ordering_timer\[23\] _1046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2933__CLK clknet_leaf_25_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3022_ _0164_ clknet_leaf_35_clock u1.ordering_timer\[18\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2806_ _0372_ _1021_ _1026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2737_ _0945_ _0983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2668_ _1206_ _0935_ _0220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1565__A2 _1163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2762__A1 _1167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1619_ u1.timer\[16\] _1237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2599_ u1.row_sel\[3\] _0877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2514__B2 spi_data_crossing\[1\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2514__A1 _0517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input39_I la_oenb[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2278__B1 _0604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2817__A2 _1025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2753__A1 _0983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2956__CLK clknet_leaf_34_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1492__B2 u1.ordering_complete\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1970_ _1197_ _0398_ _0405_ _0052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2744__A1 u1.timer\[24\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2522_ _0464_ _0826_ _0827_ spi_data_crossing\[4\].data_sync _0828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2453_ u1.ordering_complete\[24\] _0757_ _0771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2384_ _0709_ _0710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput2 io_latch_data_in net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3111__CLK clknet_leaf_29_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3005_ _0147_ clknet_leaf_35_clock u1.ordering_timer\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2432__B1 _0734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1786__A2 _1144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1594__I u0.timer_enable vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2035__I0 u1.ccr1\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2979__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1474__A1 _1096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2423__B1 _0734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2726__A1 _1321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3134__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1465__A1 _1085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1679__I u1.ccr0\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1953_ _0392_ _0393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1884_ _0311_ _0340_ _0342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2717__A1 _1303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2505_ _1041_ _0815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2436_ _1047_ _0750_ _0756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2367_ u1.ordering_complete\[13\] _0695_ _0607_ _0696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2298_ _0634_ _0635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1589__I _1206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3007__CLK clknet_leaf_4_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3157__CLK clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput191 net191 mem_write_n[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput180 net180 mem_address_right[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2644__B1 _1196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3270_ net95 net111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1922__A2 _0359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2221_ _0376_ u1.row_col_select\[9\] _0552_ _0564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2152_ _0521_ _0522_ _0523_ _0116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2083_ u0.cmd\[11\] _0478_ _0480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1438__B2 _1060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1989__A2 _0416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2985_ _0127_ clknet_leaf_19_clock u1.inverter_select\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1936_ u0.cmd\[11\] _0381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1867_ _0309_ _0328_ _0329_ _0330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput60 spi_data[28] net60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1798_ _1412_ _1414_ _0280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput71 spi_data[9] net71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2166__A2 _0530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2419_ _0741_ _0165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input21_I la_data_in[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1677__B2 _1268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output108_I net108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2652__B _1321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1601__A1 _1213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3186__D _0256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1668__A1 _1193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1668__B2 _1194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2770_ _1003_ net28 _0254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1721_ _1224_ u1.ccr0\[20\] _1338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1652_ u1.ccr1\[11\] _1269_ _1270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2788__I _1012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1583_ _1199_ u1.timer\[7\] _1200_ _1188_ _1201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_28_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3253_ u0.mem_write_n\[9\] clknet_leaf_12_clock net191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2204_ _0517_ u1.row_col_select\[1\] _0553_ _0555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3184_ _0254_ clknet_leaf_36_clock net144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2135_ u0.cmd\[15\] _0507_ _0512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2066_ u0.cmd\[6\] _0468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2084__A1 _1104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1831__A1 _0296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2968_ _0110_ clknet_leaf_28_clock u1.ordering_complete\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1919_ u0.cmd\[6\] _0369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2899_ _0041_ clknet_leaf_26_clock u1.ccr0\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input69_I spi_data[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1510__B1 u1.ordering_timer\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2822_ u0.cmd\[14\] _1017_ _1035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2862__CLK clknet_leaf_7_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2753_ _0983_ _0992_ _0993_ _0247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1704_ u1.timer\[18\] _1321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2684_ _0945_ _0946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3218__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1635_ u1.ccr1\[14\] _1253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1566_ u1.ccr1\[28\] _1173_ u1.ccr1\[24\] _1165_ _1184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3305_ net171 net181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1497_ u1.ordering_timer\[4\] _1122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_39_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3236_ u0.cmd\[18\] clknet_leaf_9_clock net164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3167_ spi_data_crossing\[24\].A clknet_leaf_10_clock spi_data_crossing\[24\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_5_clock clknet_2_0__leaf_clock clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2118_ _0474_ u1.ordering_complete\[24\] _0496_ _0502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3098_ _0232_ clknet_leaf_34_clock u1.timer\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2049_ _1133_ _0453_ _0456_ _0080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_8_clock_I clknet_2_1__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output175_I net175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2048__A1 _0454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2885__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1420_ u0.cmd\[26\] _1044_ _1045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1731__B1 u1.ccr0\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3021_ _0163_ clknet_leaf_35_clock u1.ordering_timer\[17\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2805_ _1012_ _1025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3040__CLK clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2736_ _1233_ _0980_ _0981_ _0982_ _0241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2667_ _0934_ _0935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1618_ u1.timer\[17\] _1236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2598_ u1.row_sel\[4\] _0876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3190__CLK clknet_leaf_38_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1549_ u1.timer\[30\] _1167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_45_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3219_ u1.inverter_select\[5\] clknet_leaf_21_clock net132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3063__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2126__I _0486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1965__I u0.cmd\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2744__A2 _1327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2521_ _0820_ _0827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2900__CLK clknet_leaf_25_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2452_ _0769_ _0765_ _0770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_39_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2383_ _0624_ _0709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput3 io_reset_n_in net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3004_ _0146_ clknet_leaf_34_clock u1.ordering_timer\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2680__A1 _0937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2480__B _0603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2035__I1 _0387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2719_ _0968_ _0969_ _0971_ _0235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xclkbuf_leaf_23_clock clknet_2_3__leaf_clock clknet_leaf_23_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input51_I spi_data[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_38_clock clknet_2_0__leaf_clock clknet_leaf_38_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2147__S _0514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3086__CLK clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3189__D _0259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1785__I u0.timer_enable vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2923__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2726__A2 _0282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2662__A1 u1.ccr1\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1952_ u0.cmd\[16\] _0391_ _0351_ _0392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_14_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1883_ _0330_ _0340_ _0341_ _0029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_30_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2717__A2 _0966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_35_clock_I clknet_2_0__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2504_ _0810_ _0709_ _0814_ _0177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2435_ _0624_ _0755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2350__B1 _0662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2366_ _1101_ _0685_ _0694_ _0695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2297_ _0602_ _0634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2946__CLK clknet_leaf_1_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2708__A2 _0961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput170 net170 mem_address_left[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput181 net181 mem_address_right[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput192 net192 output_active_left vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_47_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2192__I0 _0469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2644__A1 _1200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3101__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3251__CLK clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2220_ _0563_ _0144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2183__I0 _0459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2151_ _0404_ _0522_ _0523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1930__I0 u1.ccr0\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2082_ _1113_ _0453_ _0479_ _0090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_19_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2969__CLK clknet_leaf_28_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2984_ _0126_ clknet_leaf_20_clock u1.inverter_select\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2742__C _0982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1935_ _1344_ _0378_ _0380_ _0042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1866_ _1402_ _0329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput61 spi_data[29] net61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput50 spi_data[19] net50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput72 spi_data_clock net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_1797_ _1351_ u1.timer\[30\] u1.timer\[29\] _1413_ _1414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_44_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2418_ _0583_ _0719_ _0734_ _0740_ _0741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1677__A2 u1.ccr0\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2349_ _0670_ _0678_ _0679_ _0680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input14_I la_data_in[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2626__A1 u1.row_sel\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3124__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1668__A2 u1.ccr0\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1720_ _1233_ u1.ccr0\[21\] _1337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1651_ u1.timer\[11\] _1269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_28_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1582_ u1.ccr1\[6\] _1200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3252_ u0.mem_write_n\[8\] clknet_leaf_12_clock net190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2203_ _0554_ _0136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1659__A2 _1266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input6_I la_data_in[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3183_ _0253_ clknet_leaf_32_clock net146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2134_ _1078_ _0490_ _0511_ _0110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2608__B2 u1.row_sel\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2065_ _0467_ _0085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2084__A2 _0453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3147__CLK clknet_leaf_2_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2967_ _0109_ clknet_leaf_33_clock u1.ordering_complete\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2044__I _0451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1918_ _0368_ _0037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2898_ _0040_ clknet_leaf_26_clock u1.ccr0\[24\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1849_ _0311_ u1.col_limit\[5\] _0312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_11_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2147__I0 _0462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2647__C _1202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_4_clock_I clknet_2_0__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1793__I _1345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1510__A1 u1.ordering_timer\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1968__I u0.cmd\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2821_ _1301_ _1015_ _1034_ _0274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2752_ _1394_ _1345_ _1411_ _0988_ _0993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_9_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1703_ u1.ccr0\[18\] _1320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1577__B2 _1194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1577__A1 u1.ccr1\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2683_ _0933_ _0945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1634_ u1.ccr1\[15\] _1252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1565_ u1.ccr1\[25\] _1163_ _1183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3304_ net170 net180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3235_ u0.cmd\[17\] clknet_leaf_12_clock net163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1496_ u1.ordering_timer\[5\] _1121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2129__I0 _0442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3166_ net56 net72 spi_data_crossing\[24\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2039__I u0.cmd\[16\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2117_ _1054_ _0500_ _0501_ _0103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1501__B2 u1.ordering_complete\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3097_ _0231_ clknet_leaf_4_clock u1.timer\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2048_ _0454_ _0455_ _0456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1568__A1 _1183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output168_I net168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2658__B _0925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2048__A2 _0455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1731__A1 _1180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1899__S _0354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3020_ _0162_ clknet_leaf_35_clock u1.ordering_timer\[16\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2804_ _1281_ _1014_ _1024_ _0267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2750__C _0982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2735_ _0933_ _0982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2666_ _0933_ _0934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1617_ u1.ccr1\[20\] _1224_ _1232_ _1234_ _1235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_2597_ _0309_ _0874_ _1212_ _0875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1722__A1 _1237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1548_ _1165_ _1166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2478__B _0791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1479_ u1.ordering_complete\[11\] _1104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3218_ u1.inverter_select\[4\] clknet_leaf_21_clock net131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2278__A2 _0601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3149_ spi_data_crossing\[15\].A clknet_leaf_2_clock spi_data_crossing\[15\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1713__B2 u1.timer\[22\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1713__A1 _1327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2852__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3208__CLK clknet_leaf_38_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1795__A4 u1.timer\[24\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2142__I _0457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2520_ _0817_ _0826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1952__A1 u0.cmd\[16\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2451_ _1085_ _0769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_4_clock clknet_2_0__leaf_clock clknet_leaf_4_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_29_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2382_ _1059_ _0708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3003_ _0145_ clknet_leaf_23_clock u1.row_col_select\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput4 la_data_in[0] net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2680__A2 _0942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_31_clock_I clknet_2_2__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2432__A2 _0719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2718_ _0970_ _0971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1943__A1 _0385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1891__I u0.cmd\[17\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2649_ _1277_ _0916_ _0917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2875__CLK clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input44_I spi_data[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2423__A2 _0719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1934__A1 _0379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3030__CLK clknet_leaf_30_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2662__A2 _1173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2137__I _0454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3180__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1951_ u0.cmd\[17\] _0391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2414__A2 _0729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1882_ u1.col_sel\[4\] _0338_ _0341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2898__CLK clknet_leaf_26_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2503_ _0603_ _0813_ _0814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2434_ u1.ordering_timer\[22\] _0754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2365_ _0693_ _0694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2350__A1 _0675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2296_ _0633_ _0150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2102__A1 _1061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2047__I _0451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput160 net160 io_update_cycle_complete_oeb vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput171 net171 mem_address_left[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput193 net193 output_active_right vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput182 net182 mem_write_n[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__3053__CLK clknet_leaf_6_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2341__A1 _0670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1796__I u1.timer\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2832__D u1.row_sel\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2580__A1 _1160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2183__I1 u1.inverter_select\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2332__A1 _0648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2150_ _0514_ _0522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1930__I1 _0376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2081_ u0.cmd\[10\] _0478_ _0479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_22_clock clknet_2_3__leaf_clock clknet_leaf_22_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_19_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2983_ _0125_ clknet_leaf_17_clock u1.col_limit\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1934_ _0379_ _0370_ _0380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_37_clock clknet_2_0__leaf_clock clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1865_ u1.col_sel\[6\] _0310_ _0327_ _0328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput40 spi_data[0] net40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput62 spi_data[2] net62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput51 spi_data[1] net51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1796_ u1.timer\[28\] _1413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3076__CLK clknet_leaf_7_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2417_ _0735_ _0738_ _0739_ _0740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2323__A1 _1111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2348_ u1.ordering_complete\[11\] _0658_ _0679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2279_ _0618_ _0148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2913__CLK clknet_leaf_7_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2505__I _1041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_0_clock_I clknet_2_0__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2314__A1 u1.ordering_timer\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1840__A3 _0301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3099__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1650_ u1.timer\[10\] _1268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1581_ u1.ccr1\[7\] _1199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2150__I _0514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3251_ u0.mem_write_n\[7\] clknet_leaf_12_clock net189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2936__CLK clknet_leaf_28_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2202_ _0513_ u1.row_col_select\[0\] _0553_ _0554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3182_ _0252_ clknet_leaf_31_clock net148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2133_ u0.cmd\[14\] _0507_ _0511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2064_ _0466_ u1.ordering_complete\[5\] _0460_ _0467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2966_ _0108_ clknet_leaf_28_clock u1.ordering_complete\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1917_ u1.ccr0\[21\] _0367_ _0354_ _0368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2897_ _0039_ clknet_leaf_23_clock u1.ccr0\[23\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1848_ u1.col_sel\[5\] _0311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2060__I _0404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2544__B2 spi_data_crossing\[13\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2544__A1 _0385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1779_ _1350_ _1347_ _1396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2147__I1 u1.row_limit\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3241__CLK clknet_leaf_10_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2232__B1 _1111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2171__S _0529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2959__CLK clknet_leaf_33_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2820_ u0.cmd\[13\] _1029_ _1034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2751_ _1410_ _0990_ _1394_ _0992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1702_ u1.ccr0\[19\] _1319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1577__A2 _1193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2682_ _0935_ _0944_ _0225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1633_ _1247_ _1248_ _1249_ _1250_ _1251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2526__A1 _0469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1564_ _1176_ _1177_ _1179_ _1181_ _1182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__2526__B2 spi_data_crossing\[6\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3303_ net169 net179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1495_ _1108_ _1115_ _1119_ _1120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3234_ u0.cmd\[16\] clknet_leaf_8_clock net162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2129__I1 u1.ordering_complete\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3114__CLK clknet_leaf_29_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3165_ spi_data_crossing\[23\].A clknet_leaf_10_clock spi_data_crossing\[23\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2116_ u0.cmd\[7\] _0493_ _0501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3096_ _0230_ clknet_leaf_5_clock u1.timer\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2047_ _0451_ _0455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2949_ _0091_ clknet_leaf_1_clock u1.ordering_complete\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_26_clock_I clknet_2_3__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2840__D u1.col_sel\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2756__A1 _0982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3137__CLK clknet_leaf_2_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1495__A1 _1108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2803_ _0468_ _1021_ _1024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2734_ u1.timer\[21\] u1.timer\[20\] _0281_ _0976_ _0981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_30_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2665_ _1279_ _0932_ _0933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2596_ _0320_ _0872_ _0873_ _0874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1616_ u1.ccr1\[21\] _1233_ u1.ccr1\[20\] _1223_ _1234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__1970__A2 _0398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1547_ u1.timer\[24\] _1165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1478_ u1.ordering_timer\[12\] _1103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3217_ u1.inverter_select\[3\] clknet_leaf_21_clock net130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3148_ net46 net72 spi_data_crossing\[15\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1889__I u0.cmd\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3079_ _0004_ clknet_leaf_14_clock u0.run_state\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1789__A2 _1280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1477__B2 u1.ordering_complete\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2729__A1 _0281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2450_ _0768_ _0169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3254__I clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2381_ _0707_ _0161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3002_ _0144_ clknet_leaf_22_clock u1.row_col_select\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput5 la_data_in[10] net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1658__B _1274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2717_ _1303_ _0966_ _0970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_10_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2648_ _0911_ _0913_ _0915_ _0916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2489__B _0607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2579_ _0862_ _0204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input37_I la_oenb[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2508__I _0817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2431__I0 u1.ordering_complete\[21\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2726__A4 _0970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2414__A3 _0724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1950_ _1352_ _0361_ _0390_ _0047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1881_ u1.col_sel\[4\] _0338_ _0340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1925__A2 _0359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2502_ u1.ordering_complete\[31\] _0812_ _0714_ _0813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2433_ _0753_ _0167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1689__A1 _1303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1689__B2 _1254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2364_ _0676_ _1116_ _0665_ _0692_ _0693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_9_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2350__A2 _0655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1941__B _0384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2295_ _0623_ _0626_ _0604_ _0632_ _0633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2638__B1 u1.ccr1\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2102__A2 _0489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1861__A1 _0311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1861__B2 u1.col_limit\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1613__B2 _1229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2063__I _0406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2842__CLK clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput161 net161 io_update_cycle_complete_out vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput150 net150 io_driver_io_oeb[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput172 net172 mem_address_right[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_47_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput183 net183 mem_write_n[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput194 net194 row_col_select[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__2992__CLK clknet_leaf_22_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_3_clock clknet_2_0__leaf_clock clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1852__B2 u1.col_limit\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1604__A1 _1202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2080_ _0451_ _0478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1987__I _0397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2982_ _0124_ clknet_leaf_17_clock u1.col_limit\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2865__CLK clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1933_ u0.cmd\[10\] _0379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1864_ _0312_ _0325_ _0326_ _0327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput30 la_oenb[17] net30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput63 spi_data[30] net63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput52 spi_data[20] net52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1795_ _1394_ _1410_ _1411_ u1.timer\[24\] _1412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xinput41 spi_data[10] net41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2416_ u1.ordering_complete\[19\] _0687_ _0739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2347_ _0676_ _0677_ _0678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_42_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2278_ u1.ordering_timer\[2\] _0601_ _0604_ _0617_ _0618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1897__I _0352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3020__CLK clknet_leaf_35_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2011__A1 _0402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2521__I _0820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3170__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2169__S _0529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2888__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1580_ _1196_ _1190_ _1197_ u1.timer\[4\] _1198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_7_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3250_ u0.mem_write_n\[6\] clknet_leaf_12_clock net188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3262__I clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3181_ spi_data_crossing\[31\].A clknet_leaf_10_clock spi_data_crossing\[31\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2201_ _0552_ _0553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_26_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2132_ _1079_ _0500_ _0510_ _0109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2063_ _0406_ _0466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2965_ _0107_ clknet_leaf_33_clock u1.ordering_complete\[27\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3043__CLK clknet_leaf_2_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1916_ u0.cmd\[5\] _0367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2896_ _0038_ clknet_leaf_25_clock u1.ccr0\[22\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1847_ u1.col_limit\[6\] _0310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3193__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1778_ _1394_ _1343_ _1344_ _1345_ _1348_ _1395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_44_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_22_clock_I clknet_2_3__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output106_I net106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2232__B2 u1.ordering_complete\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2232__A1 _1109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_21_clock clknet_2_3__leaf_clock clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_36_clock clknet_2_0__leaf_clock clknet_leaf_36_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_48_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3066__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2471__A1 u1.ordering_complete\[26\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2750_ _1410_ _0990_ _0991_ _0982_ _0246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_13_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3257__I clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1701_ u1.timer\[19\] _1318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2681_ _1191_ _0942_ _0944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_8_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2161__I _0529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2903__CLK clknet_leaf_28_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1632_ u1.timer\[8\] _1250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1563_ u1.ccr1\[26\] _1180_ _1181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3302_ net168 net178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1494_ _1117_ _1118_ _1119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3233_ u1.row_col_select\[9\] clknet_leaf_22_clock net203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3164_ net55 net72 spi_data_crossing\[23\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2115_ _0488_ _0500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3095_ _0229_ clknet_leaf_5_clock u1.timer\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2764__C _0934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2046_ u0.cmd\[0\] _0454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2462__A1 _1085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2948_ _0090_ clknet_leaf_1_clock u1.ordering_complete\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2879_ _0013_ clknet_leaf_11_clock u0.mem_write_n\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2071__I u0.cmd\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input67_I spi_data[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2020__B _0436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3089__CLK clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2453__A1 u1.ordering_complete\[24\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2926__CLK clknet_leaf_23_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2692__A1 _0946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2802_ _1282_ _1014_ _1023_ _0266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2733_ u1.timer\[20\] _0978_ _0980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2664_ _1402_ _0927_ _0931_ _0932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2595_ _0313_ u1.col_limit\[3\] _0316_ u1.col_limit\[2\] _0315_ _0873_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1615_ _1230_ _1233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1546_ _1163_ _1164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2759__C _0934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2380__B1 _0691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3231__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1477_ _1100_ u1.ordering_complete\[14\] _1101_ u1.ordering_complete\[13\] _1102_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3216_ u1.inverter_select\[2\] clknet_leaf_22_clock net129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2267__S _0607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3147_ spi_data_crossing\[14\].A clknet_leaf_2_clock spi_data_crossing\[14\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3078_ _0006_ clknet_leaf_12_clock u0.run_state\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2066__I u0.cmd\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2029_ _1176_ _0431_ _0441_ _0075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2949__CLK clknet_leaf_1_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1789__A3 _1283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2674__A1 _0937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2851__D u0.cmd\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2729__A2 _1322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3104__CLK clknet_leaf_26_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1764__B _1380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2380_ _0703_ _0682_ _0691_ _0706_ _0707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3001_ _0143_ clknet_leaf_21_clock u1.row_col_select\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3270__I net95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2665__A1 _1279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput6 la_data_in[11] net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2417__A1 _0735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2716_ _1303_ _0966_ _0969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2647_ _1216_ _0914_ _1219_ _1202_ _0915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2578_ _0299_ _0858_ _0859_ spi_data_crossing\[26\].data_sync _0862_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_43_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1529_ u0.run_state\[4\] _1151_ _1152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2408__A1 _0711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3127__CLK clknet_leaf_38_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output98_I net98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2846__D u0.cmd\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2647__A1 _1216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_1880_ _0330_ _0338_ _0339_ _0028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_14_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2501_ _0796_ _0811_ _0805_ _0810_ _0812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2432_ u1.ordering_timer\[21\] _0719_ _0734_ _0752_ _0753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2363_ u1.ordering_timer\[13\] u1.ordering_timer\[12\] _0692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2294_ _0611_ _0628_ _0631_ _0632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1513__I u1.ordering_timer\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2638__B2 _1268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1861__A2 u1.col_limit\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2344__I u1.ordering_timer\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput151 net151 io_driver_io_oeb[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput140 net140 io_driver_io_oeb[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput195 net195 row_col_select[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput184 net184 mem_write_n[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput173 net173 mem_address_right[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput162 net162 mem_address_left[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2801__A1 _0406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_17_clock_I clknet_2_3__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2429__I _0749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2981_ _0123_ clknet_leaf_16_clock u1.col_limit\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1932_ _0358_ _0378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1863_ u1.col_sel\[6\] u1.col_limit\[6\] _0326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_37_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput20 la_data_in[8] net20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput31 la_oenb[1] net31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput64 spi_data[31] net64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput53 spi_data[21] net53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1794_ u1.timer\[25\] _1411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput42 spi_data[11] net42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2020__A2 _0430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2415_ _0736_ _0737_ _0738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_44_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2346_ _1116_ _0665_ _0677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2277_ _0611_ _0615_ _0616_ _0617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1834__A2 u0.cmd\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2074__I u0.cmd\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1598__A1 _1213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2011__A2 _0431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1522__A1 _1043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1761__A1 _1292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2200_ u0.cmd\[19\] _0485_ _0350_ _0552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_26_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3180_ net64 net72 spi_data_crossing\[31\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2131_ u0.cmd\[13\] _0507_ _0510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2062_ _0465_ _0084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2832__CLK clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1816__A2 _1144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2982__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2964_ _0106_ clknet_leaf_33_clock u1.ordering_complete\[26\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1915_ _0366_ _0036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2895_ _0037_ clknet_leaf_23_clock u1.ccr0\[21\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1846_ u1.u1.impulse_gen\[0\] _0308_ _0309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1777_ _1177_ _1394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_2_clock clknet_2_0__leaf_clock clknet_leaf_2_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1682__B _1294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2329_ _0634_ _0662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1902__S _0354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input12_I la_data_in[17] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1701__I u1.timer\[19\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1807__A2 _1409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2018__B _0435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2480__A2 _0794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2232__A2 _1110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1991__A1 _1261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1743__A1 _1167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2855__CLK clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2854__D u0.cmd\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1611__I u1.timer\[22\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2471__A2 _0757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1700_ _1299_ _1316_ _1317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2680_ _0937_ _0942_ _0943_ _0224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_8_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1631_ u1.ccr1\[8\] _1249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3301_ net167 net177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1562_ u1.timer\[26\] _1180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3273__I net104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1493_ _1111_ _1112_ _1118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3232_ u1.row_col_select\[8\] clknet_leaf_22_clock net202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3163_ spi_data_crossing\[22\].A clknet_leaf_9_clock spi_data_crossing\[22\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I la_data_in[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1498__B1 _1122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2114_ _0499_ _0102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3094_ _0228_ clknet_leaf_4_clock u1.timer\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3010__CLK clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2045_ _0452_ _0453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3160__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2947_ _0089_ clknet_leaf_0_clock u1.ordering_complete\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2352__I _0625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2878_ _0012_ clknet_leaf_11_clock u0.mem_write_n\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1973__A1 _0406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1829_ _0300_ _0302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2878__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2453__A2 _0757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2262__I _0602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2849__D u0.cmd\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3033__CLK clknet_leaf_30_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2692__A2 _0951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2437__I _0629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3183__CLK clknet_leaf_32_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2444__A2 _0750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3268__I net87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2801_ _0406_ _1021_ _1023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2732_ _0937_ _0979_ _0240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2663_ _1169_ _1172_ _1175_ _0930_ _1185_ _0931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2594_ _0322_ _0326_ _0871_ _0872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1614_ _1227_ _1231_ _1232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1707__A1 _1321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1545_ u1.timer\[25\] _1163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3215_ u1.inverter_select\[1\] clknet_leaf_20_clock net128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1476_ u1.ordering_timer\[13\] _1101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2132__A1 _1079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3146_ net45 net72 spi_data_crossing\[14\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3077_ _0218_ clknet_leaf_8_clock u0.u11.impulse_gen\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2028_ _0381_ _0423_ _0441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_20_clock clknet_2_3__leaf_clock clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_24_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1946__A1 _0387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_35_clock clknet_2_0__leaf_clock clknet_leaf_35_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output166_I net166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3056__CLK clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2123__A1 u0.cmd\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2729__A3 _0974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1937__A1 _0381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3000_ _0142_ clknet_leaf_20_clock u1.row_col_select\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput7 la_data_in[12] net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3079__CLK clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2715_ _0945_ _0968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2646_ _1210_ _1218_ _1205_ _0914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2577_ _0861_ _0203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2353__A1 _0675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1528_ _1149_ _1150_ _1151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1459_ _1075_ _1081_ _1083_ _1084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_19_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2916__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2077__I u0.cmd\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3129_ spi_data_crossing\[5\].A clknet_leaf_0_clock spi_data_crossing\[5\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2805__I _1012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2540__I _0817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_13_clock_I clknet_2_1__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2715__I _0945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3221__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2500_ u1.ordering_timer\[27\] _0783_ _0769_ _0784_ _0811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_2431_ u1.ordering_complete\[21\] _0751_ _0714_ _0752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2335__A1 _0643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2939__CLK clknet_leaf_34_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2362_ _0634_ _0691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3281__I net97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2293_ u1.ordering_complete\[4\] _0630_ _0631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2574__B2 spi_data_crossing\[24\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput130 net130 inverter_select[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_47_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2629_ _0901_ _0900_ _0902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xoutput152 net152 io_driver_io_oeb[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput141 net141 io_driver_io_oeb[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__2326__A1 _0643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput163 net163 mem_address_left[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput185 net185 mem_write_n[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput174 net174 mem_address_right[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA_input42_I spi_data[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput196 net196 row_col_select[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_29_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3244__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2801__A2 _1021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2317__A1 _0643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2857__D u0.cmd\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2980_ _0122_ clknet_leaf_17_clock u1.col_limit\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1931_ _0377_ _0041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1862_ _0315_ _0323_ _0324_ _0325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput10 la_data_in[15] net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 la_data_in[9] net21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3276__I net107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput54 spi_data[22] net54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2556__B2 spi_data_crossing\[17\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2556__A1 _0348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1793_ _1345_ _1410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput32 la_oenb[2] net32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput43 spi_data[12] net43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput65 spi_data[3] net65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2308__A1 u1.ordering_timer\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2414_ _1064_ _0729_ _0724_ _0737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__3117__CLK clknet_leaf_29_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2345_ _0675_ _0676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2276_ u1.ordering_complete\[2\] _0597_ _0616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1598__A2 _1214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2314__A4 _0627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2538__A1 _0381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2538__B2 spi_data_crossing\[11\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2130_ _0509_ _0108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2061_ _0464_ u1.ordering_complete\[4\] _0460_ _0465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2963_ _0105_ clknet_leaf_30_clock u1.ordering_complete\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1914_ u1.ccr0\[20\] _0365_ _0354_ _0366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2894_ _0036_ clknet_leaf_23_clock u1.ccr0\[20\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1845_ u1.u1.impulse_gen\[1\] _0308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1776_ _1330_ _1331_ _1342_ _1386_ _1392_ _1393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_11_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1752__A2 u1.ccr0\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2328_ _0661_ _0154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2259_ _1403_ _0595_ _0600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1807__A3 _0280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2465__B1 _0762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3121__D spi_data_crossing\[1\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1991__A2 _0416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2299__A3 _0627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2196__S _0539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1630_ u1.timer\[9\] _1248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3300_ net166 net176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1561_ _1176_ u1.timer\[27\] _1178_ u1.timer\[26\] _1179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1492_ _1116_ u1.ordering_complete\[10\] _1109_ u1.ordering_complete\[9\] _1117_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3231_ u1.row_col_select\[7\] clknet_leaf_21_clock net201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3162_ net54 net72 spi_data_crossing\[22\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2113_ _0469_ u1.ordering_complete\[22\] _0496_ _0499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3093_ _0227_ clknet_leaf_5_clock u1.timer\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2044_ _0451_ _0452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2946_ _0088_ clknet_leaf_1_clock u1.ordering_complete\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2877_ _0011_ clknet_leaf_6_clock u0.timer_enable vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1828_ _0296_ _0301_ _0013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1759_ _1363_ u1.ccr0\[1\] _1366_ _1376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1489__A1 u1.ordering_timer\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1661__A1 _1187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1964__A2 _0398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2213__I0 _0367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2972__CLK clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2718__I _0970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_1__f_clock clknet_0_clock clknet_2_1__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_1_clock clknet_2_0__leaf_clock clknet_leaf_1_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_17_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2800_ _1286_ _1014_ _1022_ _0265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2731_ _1224_ _0978_ _0979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_9_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2662_ u1.ccr1\[28\] _1173_ u1.ccr1\[27\] _1349_ _1179_ _0929_ _0930_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_8_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3284__I net100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2204__I0 _0517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2593_ _0312_ _0324_ _0870_ _0871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1613_ u1.ccr1\[23\] _1228_ u1.ccr1\[22\] _1229_ u1.ccr1\[21\] _1230_ _1231_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_1544_ _1043_ _1162_ _0007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2380__A2 _0682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3214_ u1.inverter_select\[0\] clknet_leaf_20_clock net127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1475_ u1.ordering_timer\[14\] _1100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2132__A2 _0500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3145_ spi_data_crossing\[13\].A clknet_leaf_2_clock spi_data_crossing\[13\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3076_ _0217_ clknet_leaf_7_clock u0.u11.impulse_gen\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2027_ _1178_ _0430_ _0440_ _0074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2845__CLK clknet_leaf_18_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2929_ _0071_ clknet_leaf_24_clock u1.ccr1\[23\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input72_I spi_data_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2995__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2371__A2 _0694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2123__A2 _0493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1882__A1 u1.col_sel\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3000__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3150__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput8 la_data_in[13] net8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3279__I net110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2868__CLK clknet_leaf_18_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2714_ _0958_ _0966_ _0967_ _0234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2645_ _0912_ _1198_ _1201_ _0913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2576_ u0.cmd\[25\] _0858_ _0859_ spi_data_crossing\[25\].data_sync _0861_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2353__A2 _0677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1527_ u0.run_state\[5\] _1044_ u0.run_state\[1\] _1150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1458_ u1.ordering_timer\[31\] _1073_ _1082_ _1078_ _1083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__2105__A2 _0489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3128_ net67 net72 spi_data_crossing\[5\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3059_ _0201_ clknet_leaf_9_clock u0.cmd\[23\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3023__CLK clknet_leaf_36_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2041__A1 u0.cmd\[18\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2592__A2 _0321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3173__CLK clknet_leaf_10_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2430_ _1049_ _0746_ _0750_ _0751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2361_ _0690_ _0158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2379__S _0607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2292_ _0629_ _0630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2178__I _0539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2099__A1 _0454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_34_clock clknet_2_0__leaf_clock clknet_leaf_34_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1810__I _0290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3046__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3196__CLK clknet_leaf_6_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput120 net120 data_out_right[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput131 net131 inverter_select[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2628_ u1.row_sel\[5\] _0901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput142 net142 io_driver_io_oeb[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_12_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput186 net186 mem_write_n[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput175 net175 mem_address_right[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput164 net164 mem_address_left[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2559_ _0850_ _0196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput153 net153 io_driver_io_oeb[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput197 net197 row_col_select[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input35_I la_oenb[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1876__B u1.col_sel\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1828__A1 _0296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3069__CLK clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1930_ u1.ccr0\[25\] _0376_ _0358_ _0377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2253__A1 _1212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1861_ _0311_ u1.col_limit\[5\] _0314_ u1.col_limit\[4\] _0324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2906__CLK clknet_leaf_16_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput11 la_data_in[16] net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 la_oenb[0] net22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput55 spi_data[23] net55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1792_ _1406_ _1407_ _1408_ _1409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xinput33 la_oenb[3] net33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput44 spi_data[13] net44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput66 spi_data[4] net66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3209__D _0001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2413_ u1.ordering_timer\[18\] _0723_ _0583_ _0736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2344_ u1.ordering_timer\[11\] _0675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2275_ _0612_ _0614_ _0615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3211__CLK clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2483__A1 _0796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2929__CLK clknet_leaf_24_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2235__A1 _1120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2710__A2 _0963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2060_ _0404_ _0464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2962_ _0104_ clknet_leaf_27_clock u1.ordering_complete\[24\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1913_ u0.cmd\[4\] _0365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2893_ _0035_ clknet_leaf_26_clock u1.ccr0\[19\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1844_ _0307_ net33 _0024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1775_ _1337_ _1391_ _1392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1737__B1 _1353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3234__CLK clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2327_ _0654_ _0655_ _0635_ _0660_ _0661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2258_ u1.ordering_timer\[1\] _0599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2189_ _0546_ _0130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1807__A4 _0288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2465__A1 _0774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3107__CLK clknet_leaf_24_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1431__A2 u1.ordering_complete\[20\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1560_ u1.ccr1\[26\] _1178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1491_ u1.ordering_timer\[10\] _1116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3230_ u1.row_col_select\[6\] clknet_leaf_22_clock net200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3161_ spi_data_crossing\[21\].A clknet_leaf_8_clock spi_data_crossing\[21\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2695__A1 _0946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2112_ _0498_ _0101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3092_ _0226_ clknet_leaf_5_clock u1.timer\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3222__D u1.inverter_select\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2043_ _0448_ _0450_ _0451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2447__A1 _0757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2462__A4 _0778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2945_ _0087_ clknet_leaf_2_clock u1.ordering_complete\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2876_ _0022_ clknet_leaf_9_clock u0.write_config_n vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1827_ _0299_ _1149_ _0300_ _0301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1758_ _1299_ _1316_ _1375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1689_ _1303_ _1304_ _1305_ _1254_ _1306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_1_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2686__A1 _0942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1489__A2 _1104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2438__A1 u1.ordering_complete\[22\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output104_I net104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1661__A2 _1222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2374__B1 _0691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2000__S _0423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2677__A1 _0937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1778__C _1348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2730_ _0968_ _0977_ _0978_ _0239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_9_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2661_ _0928_ _1181_ _1183_ _0929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1612_ u1.timer\[21\] _1230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2592_ u1.col_sel\[0\] _0321_ _0870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3217__D u1.inverter_select\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1543_ u0.run_state\[3\] _1144_ _1161_ _1162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1474_ _1096_ _1097_ u1.ordering_timer\[14\] _1098_ _1099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3213_ _0000_ clknet_leaf_36_clock control_trigger vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2668__A1 _1206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3144_ net44 net72 spi_data_crossing\[13\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3075_ _0216_ clknet_leaf_14_clock u1.row_sel\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2026_ _0379_ _0423_ _0440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2140__I0 _0513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2928_ _0070_ clknet_leaf_24_clock u1.ccr1\[22\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2859_ u0.cmd\[15\] clknet_leaf_19_clock net101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input65_I spi_data[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2659__A1 _1187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2198__I0 _0476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3037__D _0179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2876__D _0022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 la_data_in[14] net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1625__A2 _1237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2822__A1 u0.cmd\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2586__B1 _0865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3295__I net148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2713_ _1300_ _0963_ _1254_ _0967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2644_ _1200_ _1188_ _1196_ _1190_ _0912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2575_ _0860_ _0202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1526_ u0.cmd\[27\] _1149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1561__B2 u1.timer\[26\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1457_ u1.ordering_timer\[30\] _1082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3127_ spi_data_crossing\[4\].A clknet_leaf_38_clock spi_data_crossing\[4\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3058_ _0200_ clknet_leaf_9_clock u0.cmd\[22\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2113__I0 _0469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2009_ _0426_ _0430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2813__A1 u0.cmd\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2962__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output171_I net171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1927__I0 u1.ccr0\[24\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1552__A1 u1.ccr1\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_0_clock clknet_2_0__leaf_clock clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_8_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2568__B1 _0853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1791__A1 _1272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2360_ u1.ordering_timer\[12\] _0682_ _0662_ _0689_ _0690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2291_ _0595_ _0629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2099__A2 _0490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2835__CLK clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2985__CLK clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput110 net110 data_out_left[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_12_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1782__A1 _1171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput132 net132 inverter_select[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput121 net121 data_out_right[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_47_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2627_ _0890_ _0899_ _0900_ _0214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xoutput143 net143 io_driver_io_oeb[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput165 net165 mem_address_left[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput176 net176 mem_address_right[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_47_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2558_ u0.cmd\[18\] _0845_ _0847_ spi_data_crossing\[18\].data_sync _0850_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput154 net154 io_driver_io_oeb[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput198 net198 row_col_select[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput187 net187 mem_write_n[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2489_ _0800_ _0801_ _0607_ _0802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1509_ u1.ordering_complete\[1\] _1134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input28_I la_oenb[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3140__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output96_I net96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1773__A1 _1338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2858__CLK clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1525__A1 _1043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1828__A2 _0301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2253__A2 _0578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1860_ _0313_ u1.col_limit\[3\] _0316_ u1.col_limit\[2\] _0320_ _0322_ _0323_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_30_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 la_data_in[17] net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1791_ _1272_ _1295_ _1248_ _1250_ _1408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xinput34 la_oenb[4] net34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput23 la_oenb[10] net23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput45 spi_data[14] net45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput56 spi_data[24] net56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput67 spi_data[5] net67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2412_ _0606_ _0735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2343_ _0674_ _0156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2274_ _1136_ _0613_ _0614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3013__CLK clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3163__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1989_ _1271_ _0416_ _0417_ _0059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2827__I _1037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2483__A2 _0791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1994__A1 _0387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2794__I0 u1.ccr0\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_33_clock clknet_2_2__leaf_clock clknet_leaf_33_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1906__I u0.cmd\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3036__CLK clknet_leaf_15_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2737__I _0945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3186__CLK clknet_leaf_36_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2961_ _0103_ clknet_leaf_33_clock u1.ordering_complete\[23\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1912_ _1319_ _0359_ _0364_ _0035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2892_ _0034_ clknet_leaf_26_clock u1.ccr0\[18\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1843_ net15 _0307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1774_ _1333_ _1390_ _1391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1737__A1 _1351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1737__B2 u1.timer\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2326_ _0643_ _0657_ _0659_ _0660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2257_ _0565_ _0598_ _0146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2188_ _0365_ u1.inverter_select\[4\] _0545_ _0546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2465__A2 _0755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2382__I _1059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1976__A1 _0369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1927__S _0358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3059__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2969__D _0111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2557__I _0849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1461__I u1.ordering_complete\[24\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2292__I _0629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1967__A1 _1213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1719__A1 _1236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2392__A1 _0329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1490_ _1109_ _1110_ _1111_ _1112_ _1114_ _1115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XTAP_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3160_ net53 net72 spi_data_crossing\[21\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2467__I u1.ordering_timer\[26\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2111_ _0466_ u1.ordering_complete\[21\] _0496_ _0498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3091_ _0225_ clknet_leaf_3_clock u1.timer\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2042_ u0.write_config_n u0.cmd\[21\] u0.cmd\[20\] _0449_ _0450_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_47_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1655__B1 u1.ccr1\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3298__I net164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2944_ _0086_ clknet_leaf_2_clock u1.ordering_complete\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2875_ u0.latch_cmd clknet_leaf_8_clock u0.update_cmd vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1826_ u0.cmd\[31\] _0297_ _0300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3201__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1546__I _1163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1757_ _1317_ _1342_ _1373_ _1374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1688_ u1.ccr0\[14\] _1305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2135__A1 u0.cmd\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2919__CLK clknet_leaf_34_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2686__A2 _0947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2309_ u1.ordering_complete\[6\] _0630_ _0645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3289_ net155 net154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input10_I la_data_in[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2438__A2 _0757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1646__B1 _1261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1949__A1 _0389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2374__B2 _0701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2287__I _0624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3224__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2660_ u1.ccr1\[25\] _1164_ u1.ccr1\[24\] _1166_ _0928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_8_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1611_ u1.timer\[22\] _1229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2591_ _0869_ _0209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1542_ _1159_ _1045_ _1150_ _1160_ _1161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1473_ u1.ordering_complete\[14\] _1098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3212_ _0002_ clknet_leaf_37_clock latch_data vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2668__A2 _0935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input2_I io_latch_data_in vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3233__D u1.row_col_select\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3143_ spi_data_crossing\[12\].A clknet_leaf_2_clock spi_data_crossing\[12\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3074_ _0215_ clknet_leaf_13_clock u1.row_sel\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2025_ _0439_ _0073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2927_ _0069_ clknet_leaf_23_clock u1.ccr1\[21\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2858_ u0.cmd\[14\] clknet_leaf_19_clock net100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2789_ _0345_ _1015_ _1016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1809_ net16 net3 net34 _0290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input58_I spi_data[26] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2891__CLK clknet_leaf_25_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3247__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2283__B1 _0604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2712_ _1254_ _1300_ _1262_ _0961_ _0966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_9_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2643_ u1.ccr1\[7\] _1193_ _0911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2574_ u0.cmd\[24\] _0858_ _0859_ spi_data_crossing\[24\].data_sync _0860_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1525_ _1043_ _1148_ _0009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1561__A2 u1.timer\[27\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1456_ _1077_ _1080_ _1081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3126_ net66 net72 spi_data_crossing\[4\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3057_ _0199_ clknet_leaf_8_clock u0.cmd\[21\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__2113__I1 u1.ordering_complete\[22\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2008_ u1.ccr1\[19\] _0429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2813__A2 _1029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2390__I _0624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output164_I net164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1927__I1 _0374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2501__A1 _0796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2804__A2 _1014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2006__S _0427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1543__A2 _1144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2740__A1 _0983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2290_ _1122_ _0627_ _0628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_42_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2408__C _0716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1819__I u0.cmd\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput100 net100 data_out_left[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2626_ u1.row_sel\[4\] _0897_ _0900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_12_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1782__A2 u1.ccr0\[31\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput122 net122 data_out_right[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput111 net111 data_out_right[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput133 net133 inverter_select[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput177 net177 mem_address_right[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput166 net166 mem_address_left[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2557_ _0849_ _0195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3092__CLK clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput155 net155 io_driver_io_oeb[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput144 net144 io_driver_io_oeb[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__2031__I0 u1.ccr1\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput199 net199 row_col_select[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput188 net188 mem_write_n[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_47_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2488_ _1076_ _0796_ _1093_ _0790_ _0801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_1508_ u1.ordering_complete\[0\] _1133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1439_ u1.ordering_timer\[19\] _1064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_29_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1837__A3 _0305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2495__B1 _0805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3109_ _0243_ clknet_leaf_24_clock u1.timer\[23\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2247__B1 u1.ordering_timer\[26\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1470__A1 _1084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2722__A1 _0283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2789__A1 _0345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2253__A3 _0582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1790_ _1206_ _1208_ _1214_ _1203_ _1407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xinput13 la_data_in[1] net13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput46 spi_data[15] net46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput35 la_oenb[5] net35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput24 la_oenb[11] net24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput57 spi_data[25] net57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput68 spi_data[6] net68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2411_ _0634_ _0734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2342_ u1.ordering_timer\[10\] _0655_ _0662_ _0673_ _0674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2952__CLK clknet_leaf_35_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2273_ _1138_ _0599_ _0613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1452__B2 u1.ordering_complete\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1549__I u1.timer\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1988_ _0381_ _0413_ _0417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2609_ u1.row_sel\[6\] _0526_ _0524_ u1.row_sel\[5\] _0887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2704__A1 _1272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input40_I spi_data[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output127_I net127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1994__A2 _0394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2794__I1 _0360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2975__CLK clknet_leaf_15_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1809__I0 net16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2960_ _0102_ clknet_leaf_33_clock u1.ordering_complete\[22\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2891_ _0033_ clknet_leaf_25_clock u1.ccr0\[17\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1911_ _0363_ _0361_ _0364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1842_ _0306_ _0004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1773_ _1338_ _1389_ _1335_ _1390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1737__A2 _1352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3236__D u0.cmd\[18\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2325_ _1112_ _0658_ _0659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3130__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2256_ _1139_ _0597_ _0598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_38_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2187_ _0539_ _0545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_25_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2848__CLK clknet_leaf_23_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2998__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2464__I0 u1.ordering_complete\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1967__A2 _0398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3003__CLK clknet_leaf_23_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3153__CLK clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3090_ _0224_ clknet_leaf_5_clock u1.timer\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2110_ _0497_ _0100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2041_ u0.cmd\[18\] _0349_ _0449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2447__A3 _0765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1655__B2 _1268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2943_ _0085_ clknet_leaf_1_clock u1.ordering_complete\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2874_ _0031_ clknet_leaf_17_clock u1.col_sel\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1825_ u0.cmd\[26\] _0299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1756_ _1362_ _1372_ _1373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1687_ u1.ccr0\[15\] _1304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1562__I u1.timer\[26\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2135__A2 _0507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2308_ u1.ordering_timer\[6\] _0636_ _0644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_39_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3288_ net153 net152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2239_ _1210_ _0580_ _0581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_32_clock clknet_2_2__leaf_clock clknet_leaf_32_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3026__CLK clknet_leaf_31_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3176__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2374__A2 _0682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1472__I u1.ordering_complete\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1885__A1 _0331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2677__A3 _0941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1637__B2 _1254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2252__B _0590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1610_ u1.timer\[23\] _1228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2590_ _1040_ _0864_ _0865_ spi_data_crossing\[31\].data_sync _0869_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1541_ u0.cmd\[27\] _1160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1472_ u1.ordering_complete\[15\] _1097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3211_ _0003_ clknet_leaf_37_clock reset_n vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2117__A2 _0500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3142_ net43 net72 spi_data_crossing\[12\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3073_ _0214_ clknet_leaf_13_clock u1.row_sel\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1628__A1 _1235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2024_ u1.ccr1\[25\] _0376_ _0438_ _0439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3049__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2926_ _0068_ clknet_leaf_23_clock u1.ccr1\[20\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3199__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2857_ u0.cmd\[13\] clknet_leaf_19_clock net99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1808_ _1401_ _1403_ _0289_ _0023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_15_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2788_ _1012_ _1015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1739_ _1348_ _1350_ _1354_ _1355_ _1356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1867__A1 _0309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output207_I net207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2347__A2 _0677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2298__I _0634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2909__CLK clknet_leaf_6_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2586__A2 _0864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2711_ _0935_ _0965_ _0233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2642_ _1255_ _0909_ _1260_ _1264_ _0910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2573_ _0846_ _0859_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1524_ u0.cmd\[28\] u0.run_state\[2\] _1147_ u0.run_state\[5\] _1148_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1455_ u1.ordering_timer\[30\] _1078_ u1.ordering_timer\[29\] _1079_ _1080_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1849__A1 _0311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3125_ spi_data_crossing\[3\].A clknet_leaf_0_clock spi_data_crossing\[3\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3056_ _0198_ clknet_leaf_8_clock u0.cmd\[20\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_2007_ _0428_ _0066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2671__I _0933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2026__A1 _0379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2909_ _0051_ clknet_leaf_6_clock u1.ccr1\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input70_I spi_data[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3214__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1750__I _1214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2501__A2 _0811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2017__A1 _0369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2568__A2 _0852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1776__B1 _1342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2881__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3239__D u0.cmd\[21\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput101 net101 data_out_left[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2625_ u1.row_sel\[4\] _0897_ _0899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput112 net112 data_out_right[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput123 net123 data_out_right[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_47_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput134 net134 inverter_select[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__3237__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput167 net167 mem_address_left[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2556_ _0348_ _0845_ _0847_ spi_data_crossing\[17\].data_sync _0849_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput156 net156 io_driver_io_oeb[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput145 net145 io_driver_io_oeb[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2031__I1 _0442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput189 net189 mem_write_n[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput178 net178 mem_address_right[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__2731__A2 _0978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2487_ u1.ordering_timer\[28\] _0791_ u1.ordering_timer\[29\] _0800_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1507_ _1127_ _1130_ _1131_ _1132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1438_ u1.ordering_timer\[19\] _1058_ _1059_ _1060_ _1062_ _1063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__2495__A1 _1082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2666__I _0933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3108_ _0242_ clknet_leaf_24_clock u1.timer\[22\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3039_ _0181_ clknet_leaf_6_clock u0.cmd\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2247__A1 u1.ordering_timer\[27\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2247__B2 _0504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2486__A1 _0796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2789__A2 _1015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 la_data_in[2] net14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput36 la_oenb[6] net36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput25 la_oenb[12] net25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2410__A1 _0729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput58 spi_data[26] net58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput47 spi_data[16] net47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput69 spi_data[7] net69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2410_ _0729_ _0710_ _0733_ _0164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2013__I1 _0365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2341_ _0670_ _0671_ _0672_ _0673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2713__A2 _0963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2272_ _1138_ _0599_ u1.ordering_timer\[2\] _0612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_42_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1452__A2 u1.ordering_complete\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1987_ _0397_ _0416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2401__A1 _1068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2608_ _0524_ u1.row_sel\[5\] _0521_ u1.row_sel\[4\] _0885_ _0886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__1507__A3 _1131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2539_ _0837_ _0189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input33_I la_oenb[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2468__A1 _0774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2640__A1 _1274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1475__I u1.ordering_timer\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1682__A2 u1.ccr0\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3082__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1809__I1 net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1910_ u0.cmd\[3\] _0363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2890_ _0032_ clknet_leaf_23_clock u1.ccr0\[16\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1841_ _0304_ u0.run_state\[2\] _1155_ _0306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_30_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1772_ _1323_ _1325_ _1387_ _1388_ _1389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_38_clock_I clknet_2_0__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2324_ _0629_ _0658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2255_ _0596_ _0597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2186_ _0544_ _0129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2120__S _0488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2689__A1 u1.timer\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2942__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1933__I u0.cmd\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2040_ _0447_ _0347_ _0448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_48_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1655__A2 _1272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2604__A1 u1.row_limit\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2942_ _0084_ clknet_leaf_3_clock u1.ordering_complete\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2873_ _0030_ clknet_leaf_19_clock u1.col_sel\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2713__B _1254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1824_ _0296_ _0298_ _0012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2368__B1 _0691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1755_ _1366_ _1368_ _1371_ _1372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_11_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2004__I _0422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1686_ u1.timer\[15\] _1303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1843__I net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3287_ net151 net150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2307_ _0610_ _0643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1894__A2 u0.cmd\[18\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2238_ _1205_ _1216_ _1217_ _1220_ _0580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_26_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2143__I0 _0517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2169_ _0462_ u1.col_limit\[3\] _0529_ _0535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1646__A2 u1.timer\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2965__CLK clknet_leaf_33_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output187_I net187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1957__I0 u1.ccr1\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1637__A2 u1.timer\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2252__C _0593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3120__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1540_ u0.run_state\[6\] _1159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1471_ u1.ordering_timer\[15\] _1096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2838__CLK clknet_leaf_18_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3210_ _0279_ clknet_leaf_36_clock net137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3141_ spi_data_crossing\[11\].A clknet_leaf_2_clock spi_data_crossing\[11\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3072_ _0213_ clknet_leaf_13_clock u1.row_sel\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2988__CLK clknet_leaf_22_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2023_ _0426_ _0438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_35_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2925_ _0067_ clknet_leaf_17_clock u1.ccr1\[19\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2856_ u0.cmd\[12\] clknet_leaf_20_clock net98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1807_ _1405_ _1409_ _0280_ _0288_ _0289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_15_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2787_ _1013_ _1014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1738_ _1171_ u1.ccr0\[31\] u1.ccr0\[24\] _1166_ _1355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1669_ u1.ccr0\[4\] _1286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2816__A1 u0.cmd\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output102_I net102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_7_clock_I clknet_2_1__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3143__CLK clknet_leaf_2_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2807__A1 _1290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2283__A2 _0601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2710_ _1258_ _0963_ _0965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_12_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2641_ _1252_ _1303_ _0909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2572_ _0844_ _0858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_31_clock clknet_2_2__leaf_clock clknet_leaf_31_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1523_ control_trigger_sync\[0\] control_trigger control_trigger_sync\[1\] _1147_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1454_ u1.ordering_complete\[29\] _1079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1849__A2 u1.col_limit\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3016__CLK clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3124_ net65 net72 spi_data_crossing\[3\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3055_ _0197_ clknet_leaf_8_clock u0.cmd\[19\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_27_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3166__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2006_ u1.ccr1\[18\] _0360_ _0427_ _0428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2026__A2 _0423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2908_ _0050_ clknet_leaf_15_clock u1.ccr1\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2839_ u1.col_sel\[1\] clknet_leaf_18_clock net84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input63_I spi_data[30] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2399__I _0723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2501__A3 _0805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2017__A2 _0431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1776__B2 _1386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3039__CLK clknet_leaf_6_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3189__CLK clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1700__A1 _1299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2256__A2 _0597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1464__B1 _1088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2624_ _0890_ _0897_ _0898_ _0213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2213__S _0558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput113 net113 data_out_right[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput124 net124 data_out_right[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput102 net102 data_out_left[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_47_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1519__A1 _1070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput168 net168 mem_address_left[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput135 net135 inverter_select[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2555_ _0848_ _0194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput157 net157 io_driver_io_oeb[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput146 net146 io_driver_io_oeb[17] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput179 net179 mem_address_right[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2486_ _0796_ _0710_ _0799_ _0174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1506_ _1125_ u1.ordering_complete\[6\] _1121_ u1.ordering_complete\[5\] _1131_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__1851__I u1.col_sel\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1437_ u1.ordering_timer\[17\] _1061_ u1.ordering_timer\[16\] _1060_ _1062_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__2168__B _0534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3107_ _0241_ clknet_leaf_24_clock u1.timer\[21\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3038_ _0180_ clknet_leaf_8_clock u0.cmd\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1455__B1 u1.ordering_timer\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1758__A1 _1299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2486__A2 _0710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2238__A2 _1216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1749__A1 _1363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput15 la_data_in[3] net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 la_oenb[13] net26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput37 la_oenb[7] net37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2410__A2 _0710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1936__I u0.cmd\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput59 spi_data[27] net59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput48 spi_data[17] net48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2033__S _0438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2340_ u1.ordering_complete\[10\] _0658_ _0672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1921__A1 _0369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2767__I net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2271_ _0610_ _0611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_34_clock_I clknet_2_0__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1988__A1 _0381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3204__CLK clknet_leaf_16_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1986_ _0415_ _0058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2607_ u1.row_limit\[4\] _0876_ u1.row_limit\[3\] _0877_ _0884_ _0885_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2165__A1 _0457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2538_ _0381_ _0832_ _0833_ spi_data_crossing\[11\].data_sync _0837_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2704__A3 _0950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1581__I u1.ccr1\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2469_ _0769_ _0784_ _0785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_29_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input26_I la_oenb[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2118__S _0496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3301__I net167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1979__A1 _1199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1957__S _0394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2871__CLK clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3227__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1840_ _0304_ _1153_ _0301_ _0021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1771_ _1336_ _1334_ _1388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2323_ _1111_ _0656_ _0657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2254_ _0595_ _0596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2185_ _0363_ u1.inverter_select\[3\] _0540_ _0544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1969_ _0404_ _0400_ _0405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1576__I u1.timer\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2894__CLK clknet_leaf_23_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2689__A2 u1.timer\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2310__A1 _0643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2941_ _0083_ clknet_leaf_3_clock u1.ordering_complete\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2872_ _0029_ clknet_leaf_19_clock u1.col_sel\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1823_ u0.cmd\[31\] u0.cmd\[26\] u0.cmd\[27\] _0297_ _0298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1754_ _1364_ u1.ccr0\[0\] _1369_ _1370_ _1371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_8_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2221__S _0552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1685_ _1300_ _1301_ _1302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3286_ net149 net138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2306_ _0642_ _0151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1894__A3 u0.cmd\[21\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2237_ _1187_ _1235_ _1245_ _0579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2176__B _0538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2168_ _0319_ _0530_ _0534_ _0121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2099_ _0454_ _0490_ _0491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2690__I _0950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2359__A1 _0670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1957__I1 _0356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_3_clock_I clknet_2_0__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3072__CLK clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3173__D spi_data_crossing\[27\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2295__B1 _0604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1470_ _1084_ _1090_ _1092_ _1094_ _1095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3140_ net42 net72 spi_data_crossing\[11\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2522__B2 spi_data_crossing\[4\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2522__A1 _0464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2775__I net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3071_ _0212_ clknet_leaf_13_clock u1.row_sel\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2022_ _0437_ _0072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2825__A2 _1015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2924_ _0066_ clknet_leaf_26_clock u1.ccr1\[18\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2855_ u0.cmd\[11\] clknet_leaf_19_clock net97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1806_ _0284_ _0287_ _0288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2786_ _1012_ _1013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2061__I0 _0464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1854__I u1.col_sel\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3095__CLK clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2761__A1 u1.timer\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1737_ _1351_ _1352_ _1353_ u1.timer\[30\] _1354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1668_ _1193_ u1.ccr0\[7\] u1.ccr0\[4\] _1194_ _1284_ _1285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1599_ _1207_ u1.ccr1\[0\] _1217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3269_ net88 net94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2932__CLK clknet_leaf_25_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2816__A2 _1029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2752__A1 _1394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2796__S _1013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2807__A2 _1025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2268__B1 _0604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1939__I _0353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2440__B1 _0734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2640_ _1274_ _1251_ _1275_ _0907_ _0908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2571_ _0857_ _0201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1522_ _1043_ _1146_ _0010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1453_ u1.ordering_complete\[30\] _1078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2955__CLK clknet_leaf_33_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3123_ spi_data_crossing\[2\].A clknet_leaf_38_clock spi_data_crossing\[2\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3054_ _0196_ clknet_leaf_8_clock u0.cmd\[18\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2005_ _0426_ _0427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_35_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2907_ _0049_ clknet_leaf_15_clock u1.ccr1\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2838_ u1.col_sel\[0\] clknet_leaf_18_clock net83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2769_ net10 _1003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input56_I spi_data[24] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_29_clock_I clknet_2_2__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3304__I net170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3110__CLK clknet_leaf_24_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output212_I net212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2978__CLK clknet_leaf_18_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1528__A2 _1150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2725__A1 _1322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1464__B2 u1.ordering_complete\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1767__A2 _1308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2623_ u1.row_sel\[3\] _0895_ _0898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput114 net114 data_out_right[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput125 net125 data_out_right[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput103 net103 data_out_left[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2554_ _0447_ _0845_ _0847_ spi_data_crossing\[16\].data_sync _0848_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1519__A2 _1095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2716__A1 _1303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput136 net136 inverter_select[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput158 net158 io_latch_data_oeb vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput147 net147 io_driver_io_oeb[18] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_1505_ _1128_ u1.ordering_complete\[3\] _1122_ u1.ordering_complete\[4\] _1129_ _1130_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xoutput169 net169 mem_address_left[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA_clkbuf_leaf_30_clock_I clknet_2_2__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2485_ u1.ordering_complete\[28\] _0720_ _0603_ _0798_ _0799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3133__CLK clknet_leaf_2_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1436_ u1.ordering_complete\[17\] _1061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_29_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3106_ _0240_ clknet_leaf_24_clock u1.timer\[20\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3037_ _0179_ clknet_leaf_15_clock u0.cmd\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1455__B2 _1079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output162_I net162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_30_clock clknet_2_2__leaf_clock clknet_leaf_30_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_15_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1997__A2 _0400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3006__CLK clknet_leaf_4_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput16 la_data_in[4] net16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput27 la_oenb[14] net27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput49 spi_data[18] net49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput38 la_oenb[8] net38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3156__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2270_ _0596_ _0610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1437__B2 _1060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1988__A2 _0413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1985_ u1.ccr1\[10\] _0379_ _0397_ _0415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2606_ _0880_ _0882_ _0883_ _0884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2023__I _0426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2537_ _0836_ _0188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1912__A2 _0359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2468_ _0774_ _0761_ u1.ordering_timer\[22\] _0749_ _0784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1419_ control_trigger_sync\[0\] control_trigger control_trigger_sync\[1\] _1044_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_29_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2399_ _0723_ _0724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input19_I la_data_in[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1428__B2 u1.ordering_complete\[21\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1428__A1 _1047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3029__CLK clknet_leaf_30_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3179__CLK clknet_leaf_10_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1600__A1 u1.ccr1\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output87_I net87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2459__A3 _0775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1667__B2 _1283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1667__A1 _1280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2219__I0 _0374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1770_ _1323_ _1326_ _1387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2322_ _0648_ _0649_ _0656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2253_ _1212_ _0578_ _0582_ _0594_ _0595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2184_ _0543_ _0128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1658__A1 u1.ccr1\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2219__S _0552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2607__B1 u1.row_limit\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2083__A1 u0.cmd\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1968_ u0.cmd\[4\] _0404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1899_ u1.ccr0\[16\] _0345_ _0354_ _0355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2138__A2 _0348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2689__A3 _0941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2129__S _0488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2377__A2 _0694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2598__I u1.row_sel\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1888__A1 _0331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2940_ _0082_ clknet_leaf_4_clock u1.ordering_complete\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2871_ _0028_ clknet_leaf_19_clock u1.col_sel\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1822_ _0295_ u0.update_cmd _0297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2368__A2 _0682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1753_ _1204_ u1.ccr0\[2\] _1370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1684_ u1.ccr0\[13\] _1301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2502__S _0714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3285_ net101 net117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2305_ u1.ordering_timer\[5\] _0626_ _0635_ _0641_ _0642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1894__A4 u0.cmd\[20\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2236_ _0566_ _0577_ _0578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_26_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2167_ _0399_ _0531_ _0534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2098_ _0487_ _0490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2861__CLK clknet_leaf_2_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3217__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1960__I _0397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3070_ _0211_ clknet_leaf_13_clock u1.row_sel\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1730__B1 u1.ccr0\[24\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2021_ u1.ccr1\[24\] _0374_ _0427_ _0437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2791__I _1012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2884__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2923_ _0065_ clknet_leaf_17_clock u1.ccr1\[17\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2854_ u0.cmd\[10\] clknet_leaf_19_clock net96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1805_ _0285_ _0286_ u1.timer\[21\] u1.timer\[20\] _0287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_2785_ _1011_ _1012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1736_ u1.ccr0\[30\] _1353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1667_ _1280_ _1281_ _1282_ _1283_ _1284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_28_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1598_ _1213_ _1214_ _1215_ _1203_ _1216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3268_ net87 net93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2219_ _0374_ u1.row_col_select\[8\] _0552_ _0563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3199_ _0269_ clknet_leaf_27_clock u1.ccr0\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2277__A1 _0611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_25_clock_I clknet_2_3__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output192_I net192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2650__B _0910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2752__A2 _1345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3184__D _0254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2504__A2 _0709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2570_ u0.cmd\[23\] _0852_ _0853_ spi_data_crossing\[23\].data_sync _0857_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1521_ u0.run_state\[6\] _1045_ _1145_ u0.run_state\[3\] _1146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1452_ _1076_ u1.ordering_complete\[29\] _1071_ u1.ordering_complete\[28\] _1077_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2786__I _1012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3122_ net62 net72 spi_data_crossing\[2\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3053_ _0195_ clknet_leaf_6_clock u0.cmd\[17\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2259__A1 _1403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2004_ _0422_ _0426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1482__A2 u1.ordering_complete\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3062__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2906_ _0048_ clknet_leaf_16_clock u1.ccr1\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2837_ u1.row_sel\[5\] clknet_leaf_13_clock net209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2768_ _1002_ net29 _0253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1719_ _1236_ u1.ccr0\[17\] _1336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2699_ _0946_ _0956_ _0957_ _0229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_input49_I spi_data[18] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2498__A1 _0565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2670__A1 _0935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2422__A1 _0735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2725__A2 _0974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3085__CLK clknet_leaf_38_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2661__A1 _0928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1464__A2 u1.ordering_complete\[26\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2622_ u1.row_sel\[3\] _0895_ _0897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2922__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput104 net104 data_out_left[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput115 net115 data_out_right[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2553_ _0846_ _0847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1519__A3 _1120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2716__A2 _0966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput126 net126 data_out_right[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput137 net137 io_control_trigger_oeb vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput159 net159 io_reset_n_oeb vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput148 net148 io_driver_io_oeb[19] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_1504_ _1124_ u1.ordering_complete\[7\] _1129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2484_ _0597_ _0797_ _0798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1435_ u1.ordering_complete\[16\] _1060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_3105_ _0239_ clknet_leaf_26_clock u1.timer\[19\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3036_ _0178_ clknet_leaf_15_clock u0.cmd\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2652__A1 _0429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2707__A2 _0961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2643__A1 u1.ccr1\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2945__CLK clknet_leaf_2_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput17 la_data_in[5] net17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 la_oenb[15] net28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput39 la_oenb[9] net39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1438__C _1062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1437__A2 _1061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1984_ _1247_ _0409_ _0414_ _0057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2605_ u1.row_limit\[3\] _0877_ u1.row_limit\[2\] _0881_ _0883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3100__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2536_ _0379_ _0832_ _0833_ spi_data_crossing\[10\].data_sync _0836_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3250__CLK clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2570__B1 _0853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2467_ u1.ordering_timer\[26\] _0783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1418_ _1040_ u0.cmd\[30\] _1042_ _1043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_29_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2173__I0 _0466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2468__A4 _0749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2398_ _1096_ u1.ordering_timer\[14\] _0693_ _0722_ _0723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_29_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2625__A1 u1.row_sel\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3019_ _0161_ clknet_leaf_35_clock u1.ordering_timer\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1428__A2 u1.ordering_complete\[22\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2968__CLK clknet_leaf_28_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2459__A4 _0692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2616__A1 _0891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1419__A2 control_trigger vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2092__A2 _0455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2219__I1 u1.row_col_select\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3123__CLK clknet_leaf_38_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2321_ _0625_ _0655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2252_ _1095_ _0588_ _0590_ _0593_ _0594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2183_ _0459_ u1.inverter_select\[2\] _0540_ _0543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1658__A2 _1267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2743__B u1.timer\[24\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2083__A2 _0478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1967_ _1213_ _0398_ _0403_ _0051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2386__A3 _0694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1898_ _0353_ _0354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2519_ _0825_ _0181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2689__A4 _0947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input31_I la_oenb[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3146__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1821__A2 u0.cmd\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2145__S _0514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3187__D _0257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2870_ _0027_ clknet_leaf_19_clock u1.col_sel\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2055__S _0460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1821_ u0.cmd\[28\] u0.cmd\[29\] _0296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3097__D _0231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1752_ _1367_ u1.ccr0\[3\] _1369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1683_ u1.timer\[13\] _1300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3019__CLK clknet_leaf_35_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3284_ net100 net116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2304_ _0611_ _0639_ _0640_ _0641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2828__A1 net13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2235_ _1120_ _0570_ _0573_ _0576_ _0577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3169__CLK clknet_leaf_10_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2166_ _0318_ _0530_ _0533_ _0120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2097_ _0488_ _0489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1868__I _0330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2999_ _0141_ clknet_leaf_22_clock u1.row_col_select\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1567__A1 u1.ccr1\[31\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2367__I0 u1.ordering_complete\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_21_clock_I clknet_2_3__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2648__B _0915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2819__A1 _1310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2020_ _1225_ _0430_ _0436_ _0071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2922_ _0064_ clknet_leaf_17_clock u1.ccr1\[16\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1797__A1 _1351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2853_ u0.cmd\[9\] clknet_leaf_17_clock net110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2784_ _0447_ _0347_ _0351_ _1011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1804_ u1.timer\[22\] _0286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1735_ u1.ccr0\[31\] _1352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2312__I _0647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1666_ _1190_ _1283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1597_ u1.ccr1\[2\] _1215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3267_ net86 net92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2218_ _0562_ _0143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3198_ _0268_ clknet_leaf_6_clock u1.ccr0\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2149_ u1.row_limit\[4\] _0521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2029__A2 _0431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2268__A2 _0601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2440__A2 _0755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1520_ _1144_ _1145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1971__I u0.cmd\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1451_ u1.ordering_timer\[29\] _1076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3121_ spi_data_crossing\[1\].A clknet_leaf_0_clock spi_data_crossing\[1\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2851__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3052_ _0194_ clknet_leaf_8_clock u0.cmd\[16\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2003_ _0425_ _0065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3207__CLK clknet_leaf_38_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2307__I _0610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2905_ _0047_ clknet_leaf_27_clock u1.ccr0\[31\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2751__B _1394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2836_ u1.row_sel\[4\] clknet_leaf_13_clock net208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2767_ net11 _1002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1718_ _1233_ u1.ccr0\[21\] u1.ccr0\[20\] _1224_ _1335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2734__A3 _0281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2698_ _1248_ _0954_ _0957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1649_ u1.timer\[8\] _1267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2498__A2 _0601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1458__B1 _1082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output100_I net100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2874__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2413__A2 _0723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2621_ _0890_ _0895_ _0896_ _0212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2177__A1 u0.cmd\[19\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput116 net116 data_out_right[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput105 net105 data_out_left[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2552_ _0819_ _0846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput127 net127 inverter_select[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_49_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1924__A1 _0372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput149 net149 io_driver_io_oeb[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput138 net138 io_driver_io_oeb[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_12_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1503_ u1.ordering_timer\[3\] _1128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2483_ _0796_ _0791_ _0797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1434_ u1.ordering_timer\[16\] _1059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3104_ _0238_ clknet_leaf_26_clock u1.timer\[18\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3035_ _0177_ clknet_leaf_30_clock u1.ordering_timer\[31\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2101__A1 _0457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2819_ _1310_ _1025_ _1033_ _0273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input61_I spi_data[29] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2897__CLK clknet_leaf_23_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output148_I net148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2656__B _1227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2643__A2 _1193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput18 la_data_in[6] net18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput29 la_oenb[16] net29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2159__A1 _0447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3052__CLK clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2331__A1 _1109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2058__S _0460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2398__A1 _1096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1983_ u0.cmd\[9\] _0413_ _0414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2604_ u1.row_limit\[2\] _0881_ u1.row_limit\[1\] _0878_ _0882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2535_ _0835_ _0187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2466_ _0782_ _0171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1417_ _1041_ _1042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2173__I1 u1.col_limit\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2322__A1 _0648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2397_ _1068_ _1059_ _0722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3018_ _0160_ clknet_leaf_35_clock u1.ordering_timer\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2431__S _0714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3075__CLK clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2912__CLK clknet_leaf_7_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_16_clock_I clknet_2_2__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2320_ u1.ordering_timer\[8\] _0654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2251_ _1083_ _0592_ _1074_ _0593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2304__A1 _0611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2182_ _0542_ _0127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1902__I1 _0356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1966_ _0402_ _0400_ _0403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1897_ _0352_ _0353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3098__CLK clknet_leaf_34_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2050__I u0.cmd\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2518_ _0462_ _0818_ _0821_ spi_data_crossing\[3\].data_sync _0825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2449_ _0761_ _0755_ _0762_ _0767_ _0768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2935__CLK clknet_leaf_28_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input24_I la_oenb[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2782__A1 _1009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2534__A1 _0476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3240__CLK clknet_leaf_10_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1820_ _1040_ _0295_ u0.update_cmd _0022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1751_ _1367_ u1.ccr0\[3\] u1.ccr0\[2\] _1204_ _1368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_7_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1682_ _1293_ u1.ccr0\[9\] _1294_ _1298_ _1299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2958__CLK clknet_leaf_34_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2303_ u1.ordering_complete\[5\] _0630_ _0640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3283_ net99 net115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2234_ _1114_ _0575_ _1108_ _0576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2165_ _0457_ _0531_ _0533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2096_ _0487_ _0488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2998_ _0140_ clknet_leaf_21_clock u1.row_col_select\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2064__I0 _0466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1567__A2 _1171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1949_ _0389_ _0383_ _0390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2764__A1 _1351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1811__I0 net17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2516__A1 _0459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2516__B2 spi_data_crossing\[2\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2819__A2 _1025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3113__CLK clknet_leaf_24_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1794__I u1.timer\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2055__I0 _0459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1730__A2 u1.ccr0\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2921_ _0063_ clknet_leaf_27_clock u1.ccr1\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1797__A2 u1.timer\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2852_ u0.cmd\[8\] clknet_leaf_20_clock net109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2783_ u1.ccr0\[0\] _1010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1803_ _1327_ _0285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1734_ u1.timer\[31\] _1351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1665_ u1.ccr0\[5\] _1282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1596_ u1.timer\[3\] _1214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3136__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3266_ net85 net91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2217_ _0472_ u1.row_col_select\[7\] _0558_ _0562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3197_ _0267_ clknet_leaf_15_clock u1.ccr0\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2148_ _0520_ _0115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2079_ _0477_ _0089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2037__I0 u1.ccr1\[31\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3009__CLK clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2728__A1 _0281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3159__CLK clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1450_ _1071_ u1.ordering_complete\[28\] _1072_ u1.ordering_complete\[27\] _1074_
+ _1075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_3120_ net51 net72 spi_data_crossing\[1\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3051_ _0193_ clknet_leaf_3_clock u0.cmd\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2002_ u1.ccr1\[17\] _0356_ _0423_ _0425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1467__A1 _1088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2904_ _0046_ clknet_leaf_28_clock u1.ccr0\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2835_ u1.row_sel\[3\] clknet_leaf_13_clock net207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2719__A1 _0968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2766_ _1001_ net30 _0252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1717_ _1236_ u1.ccr0\[17\] u1.ccr0\[16\] _1237_ _1334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2734__A4 _0976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2697_ _0951_ _0955_ _0956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1648_ _1260_ _1265_ _1266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1579_ u1.ccr1\[4\] _1197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2498__A3 _0808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3249_ u0.mem_write_n\[5\] clknet_leaf_13_clock net187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1458__A1 u1.ordering_timer\[31\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1697__A1 _1267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1449__A1 u1.ordering_timer\[31\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2661__A3 _1183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2620_ u1.row_sel\[1\] _0892_ u1.row_sel\[2\] _0896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput106 net106 data_out_left[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2551_ _0844_ _0845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1982__I _0393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput117 net117 data_out_right[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput128 net128 inverter_select[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput139 net139 io_driver_io_oeb[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_1502_ _1123_ _1126_ _1127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2482_ _1071_ _0796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1433_ u1.ordering_complete\[19\] _1058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3103_ _0237_ clknet_leaf_27_clock u1.timer\[17\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3034_ _0176_ clknet_leaf_33_clock u1.ordering_timer\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2101__A2 _0490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2053__I _0399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2818_ u0.cmd\[12\] _1029_ _1033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2168__A2 _0530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2749_ _1410_ _0990_ _0991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input54_I spi_data[22] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2340__A2 _0658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1603__A1 _1212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2391__C _0716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput19 la_data_in[7] net19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2841__CLK clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2159__A2 _0348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2991__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_12_clock_I clknet_2_1__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2398__A2 u1.ordering_timer\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1982_ _0393_ _0413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2603_ u1.row_sel\[2\] _0881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2601__I u1.row_sel\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2534_ _0476_ _0832_ _0833_ spi_data_crossing\[9\].data_sync _0835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2570__A2 _0852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2465_ _0774_ _0755_ _0762_ _0781_ _0782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1416_ reset_n_sync\[1\] reset_n_sync\[0\] reset_n _1041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2396_ _0708_ _0712_ _0721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3017_ _0159_ clknet_leaf_37_clock u1.ordering_timer\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2389__A2 _0714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2864__CLK clknet_leaf_15_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2511__I _0820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1824__A1 _0296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2250_ _1077_ _0591_ _0592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2069__S _0470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2181_ _0517_ u1.inverter_select\[1\] _0540_ _0542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2887__CLK clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1815__A1 net19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1500__I u1.ordering_timer\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1965_ u0.cmd\[3\] _0402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2240__A1 _1202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1896_ _0346_ _0348_ _0351_ _0352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2517_ _0824_ _0180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1751__B1 u1.ccr0\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2448_ _1054_ _0720_ _0766_ _0767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2487__B u1.ordering_timer\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2379_ u1.ordering_complete\[15\] _0705_ _0607_ _0706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input17_I la_data_in[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3042__CLK clknet_leaf_7_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3192__CLK clknet_leaf_16_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1750_ _1214_ _1367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1681_ _1295_ _1296_ _1297_ _1298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2302_ _0636_ _0638_ _0639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3282_ net98 net114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I la_data_in[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2233_ _1117_ _0574_ _0575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2289__A1 u1.ordering_timer\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2164_ _0321_ _0530_ _0532_ _0119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2095_ _0486_ _0487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3065__CLK clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2997_ _0139_ clknet_leaf_20_clock u1.row_col_select\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1948_ u0.cmd\[15\] _0389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1879_ u1.col_sel\[3\] _0336_ _0339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1811__I1 net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2902__CLK clknet_leaf_29_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2452__A1 _0769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3088__CLK clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2920_ _0062_ clknet_leaf_33_clock u1.ccr1\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1797__A3 u1.timer\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2851_ u0.cmd\[7\] clknet_leaf_17_clock net108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2925__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1802_ _0281_ _1322_ _0282_ _0283_ _0284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_2782_ _1009_ net39 _0260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1733_ _1173_ u1.ccr0\[28\] u1.ccr0\[27\] _1349_ _1350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2810__S _1013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1664_ u1.ccr0\[6\] _1281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1595_ u1.ccr1\[3\] _1213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3265_ net84 net90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2216_ _0561_ _0142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3196_ _0266_ clknet_leaf_6_clock u1.ccr0\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2147_ _0462_ u1.row_limit\[3\] _0514_ _0520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2682__A1 _0935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2078_ _0476_ _1110_ _0470_ _0477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2037__I1 _0389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3230__CLK clknet_leaf_22_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2673__A1 _1206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2948__CLK clknet_leaf_1_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2728__A2 _0976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3050_ _0192_ clknet_leaf_4_clock u0.cmd\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2001_ _0424_ _0064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3260__I clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2664__A1 _1402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1467__A2 u1.ordering_complete\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2903_ _0045_ clknet_leaf_28_clock u1.ccr0\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2834_ u1.row_sel\[2\] clknet_leaf_13_clock net206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3103__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2765_ net12 _1001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1716_ _1330_ _1332_ _1333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2696_ _1293_ _1267_ _0955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3253__CLK clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1647_ _1261_ _1262_ _1264_ _1265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1578_ u1.ccr1\[5\] _1196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3248_ u0.mem_write_n\[4\] clknet_leaf_13_clock net186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3179_ spi_data_crossing\[30\].A clknet_leaf_10_clock spi_data_crossing\[30\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1458__A2 _1073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output190_I net190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2194__I0 _0472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1697__A2 u1.ccr0\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2836__D u1.row_sel\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1449__A2 _1073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3126__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1621__A2 u1.timer\[19\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput107 net107 data_out_left[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2550_ _0816_ _0844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput129 net129 inverter_select[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput118 net118 data_out_right[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__3255__I clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2481_ _1093_ _0710_ _0795_ _0173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1501_ _1124_ u1.ordering_complete\[7\] _1125_ u1.ordering_complete\[6\] _1126_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1432_ _1052_ _1053_ _1056_ _1057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__2185__I0 _0363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3102_ _0236_ clknet_leaf_27_clock u1.timer\[16\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2637__A1 _0905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3033_ _0175_ clknet_leaf_30_clock u1.ordering_timer\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2762__C _0934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2817_ _1031_ _1025_ _1032_ _0272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2748_ _0983_ _0989_ _0990_ _0245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_11_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2679_ _1287_ _0941_ _0943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input47_I spi_data[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3149__CLK clknet_leaf_2_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1603__A2 _1216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2564__B1 _0853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1981_ _1249_ _0409_ _0412_ _0056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2398__A3 _0693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2602_ u1.row_limit\[1\] _0878_ u1.row_limit\[0\] _0879_ _0880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_6_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2533_ _0834_ _0186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2464_ u1.ordering_complete\[25\] _0780_ _0714_ _0781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1415_ u0.cmd\[31\] _1040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2395_ _0610_ _0720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1530__A1 _1043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2329__I _0634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3016_ _0158_ clknet_leaf_37_clock u1.ordering_timer\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3100__D _0234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1824__A2 _0298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2180_ _0541_ _0126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1512__A1 _1128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1964_ _1215_ _0398_ _0401_ _0050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2240__A2 _1277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1895_ _0349_ _0350_ _0351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2379__I0 u1.ordering_complete\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2516_ _0459_ _0818_ _0821_ spi_data_crossing\[2\].data_sync _0824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1751__B2 _1204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2447_ _0757_ _0764_ _0765_ _0766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_25_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2378_ _0703_ _0704_ _0705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1898__I _0353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1806__A2 _0287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2981__CLK clknet_leaf_16_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2231__A2 u1.ordering_complete\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1990__A1 u0.cmd\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1742__A1 u1.timer\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1742__B2 u1.timer\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2844__D u0.cmd\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1981__A1 _1249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1680_ _1269_ u1.ccr0\[11\] _1297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2301_ _1121_ _0637_ _0638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1733__A1 _1173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3281_ net97 net113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3263__I clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2854__CLK clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2232_ _1109_ _1110_ _1111_ u1.ordering_complete\[8\] _0574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2289__A2 u1.ordering_timer\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2163_ _0454_ _0531_ _0532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2808__S _1013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2094_ _0485_ _0450_ _0486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2461__A2 _0729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2996_ _0138_ clknet_leaf_20_clock u1.row_col_select\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1947_ _1353_ _0361_ _0388_ _0046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1878_ u1.col_sel\[3\] _0336_ _0338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_31_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2452__A2 _0765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1963__A1 _0399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2839__D u1.col_sel\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2877__CLK clknet_leaf_6_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1715__A1 _1229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2427__I _0747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2850_ u0.cmd\[6\] clknet_leaf_20_clock net107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1801_ u1.timer\[16\] _0283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3258__I clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2162__I _0528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2781_ net21 _1009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1732_ _1177_ _1349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1663_ _1188_ _1280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1594_ u0.timer_enable _1212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1706__B2 _1322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3264_ net83 net89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2215_ _0369_ u1.row_col_select\[6\] _0558_ _0561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3032__CLK clknet_leaf_30_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3195_ _0265_ clknet_leaf_6_clock u1.ccr0\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2131__A1 u0.cmd\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2146_ _0519_ _0114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2077_ u0.cmd\[9\] _0476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3182__CLK clknet_leaf_31_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2979_ _0121_ clknet_leaf_17_clock u1.col_limit\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2425__A2 _0737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1633__B1 _1249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3055__CLK clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2000_ u1.ccr1\[16\] _0345_ _0423_ _0424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2416__A2 _0687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2902_ _0044_ clknet_leaf_29_clock u1.ccr0\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2833_ u1.row_sel\[1\] clknet_leaf_13_clock net205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2764_ _1351_ _0999_ _1000_ _0934_ _0251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1715_ _1229_ u1.ccr0\[22\] _1331_ _1332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2695_ _0946_ _0953_ _0954_ _0228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1646_ _1263_ u1.timer\[13\] _1261_ u1.timer\[12\] _1264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1577_ u1.ccr1\[7\] _1193_ u1.ccr1\[4\] _1194_ _1195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3247_ u0.mem_write_n\[3\] clknet_leaf_11_clock net185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2495__C _0725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2104__A1 _0399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3178_ net63 net72 spi_data_crossing\[30\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2067__I _0468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2129_ _0442_ u1.ordering_complete\[28\] _0488_ _0509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2407__A2 _0725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3078__CLK clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2530__I _0817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2915__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2852__D u0.cmd\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput119 net119 data_out_right[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput108 net108 data_out_left[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2480_ _0793_ _0794_ _0603_ _0795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1500_ u1.ordering_timer\[6\] _1125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1431_ _1050_ u1.ordering_complete\[20\] _1055_ _1056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2185__I1 u1.inverter_select\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2334__A1 _1110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput90 net90 col_select_right[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_3101_ _0235_ clknet_leaf_27_clock u1.timer\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3271__I net102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3032_ _0174_ clknet_leaf_30_clock u1.ordering_timer\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3220__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2816_ u0.cmd\[11\] _1029_ _1032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2747_ _1411_ _0988_ _0990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2678_ _1287_ _0941_ _0942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1629_ u1.ccr1\[9\] _1247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2325__A1 _1112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2938__CLK clknet_leaf_34_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2800__A2 _1014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2564__A1 u0.cmd\[20\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2847__D u0.cmd\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1914__I1 _0365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3243__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1980_ u0.cmd\[8\] _0407_ _0412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2435__I _0624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2601_ u1.row_sel\[0\] _0879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2532_ _0474_ _0832_ _0833_ spi_data_crossing\[8\].data_sync _0834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2463_ _0774_ _0779_ _0780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2394_ _0625_ _0719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1514__I _1138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3015_ _0157_ clknet_leaf_37_clock u1.ordering_timer\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2345__I _0675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2080__I _0451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2546__B2 spi_data_crossing\[14\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2546__A1 _0387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3116__CLK clknet_leaf_29_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output146_I net146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2085__I0 _0442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1512__A2 u1.ordering_complete\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2473__B1 _0762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1963_ _0399_ _0400_ _0401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1894_ u0.write_config_n u0.cmd\[18\] u0.cmd\[21\] u0.cmd\[20\] _0350_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_18_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2240__A3 _0579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2528__A1 _0472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2528__B2 spi_data_crossing\[7\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3139__CLK clknet_leaf_2_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2515_ _0823_ _0179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1751__A2 u1.ccr0\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2446_ _0761_ _0754_ _0750_ _0765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_29_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_2_0__f_clock clknet_0_clock clknet_2_0__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2377_ _0698_ _0694_ _0704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1990__A2 _0413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2455__B1 _0762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2058__I0 _0462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1773__B _1335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3280_ net96 net112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2300_ _0623_ _0627_ _0637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2231_ _0571_ u1.ordering_complete\[15\] _1099_ _0572_ _0573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2162_ _0528_ _0531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1999__I _0422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2093_ _0346_ _0347_ _0485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_4_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2461__A3 _0777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2995_ _0137_ clknet_leaf_21_clock u1.row_col_select\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1946_ _0387_ _0383_ _0388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1877_ _0330_ _0336_ _0337_ _0027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2221__I0 _0376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2429_ _0749_ _0750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input22_I la_oenb[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output109_I net109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1963__A2 _0400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_2_3__f_clock_I clknet_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1813__S net36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2855__D u0.cmd\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1800_ u1.timer\[17\] _0282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2443__I _0602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2780_ _1008_ net23 _0259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1731_ _1180_ u1.ccr0\[26\] u1.ccr0\[25\] _1164_ _1348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_15_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1662_ _1279_ u1.ccr1_flag vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3274__I net105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1593_ _1205_ _1210_ _1211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3263_ clknet_leaf_12_clock net82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2214_ _0560_ _0141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2971__CLK clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3194_ _0264_ clknet_leaf_16_clock u1.ccr0\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2145_ _0459_ u1.row_limit\[2\] _0514_ _0519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2131__A2 _0507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2076_ _0475_ _0088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2978_ _0120_ clknet_leaf_18_clock u1.col_limit\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1929_ u0.cmd\[9\] _0376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1881__A1 u1.col_sel\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2464__S _0714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1633__A1 _1247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2263__I _0603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2844__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2994__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2664__A3 _0931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1872__A1 _0331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2901_ _0043_ clknet_leaf_29_clock u1.ccr0\[27\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3269__I net88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2832_ u1.row_sel\[0\] clknet_leaf_13_clock net204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2763_ _1351_ _0999_ _1000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1714_ _1327_ _1328_ _1331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2694_ _1250_ _0951_ _0954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1645_ u1.ccr1\[13\] _1263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1576_ u1.timer\[4\] _1194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3246_ u0.mem_write_n\[2\] clknet_leaf_11_clock net184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2104__A2 _0493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3177_ spi_data_crossing\[29\].A clknet_leaf_12_clock spi_data_crossing\[29\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2128_ _0506_ _0500_ _0508_ _0107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_2059_ _0463_ _0083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2867__CLK clknet_leaf_38_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2040__A1 _0447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1551__B1 u1.ccr1\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2258__I u1.ordering_timer\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1909__A2 _0359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3022__CLK clknet_leaf_35_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput109 net109 data_out_left[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__3172__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1430_ u1.ordering_timer\[23\] _1054_ _1055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2334__A2 _0658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput80 net80 clock_out[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput91 net91 col_select_right[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__1542__B1 _1150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3100_ _0234_ clknet_leaf_27_clock u1.timer\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3031_ _0173_ clknet_leaf_30_clock u1.ordering_timer\[27\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2815_ u1.ccr0\[11\] _1031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2746_ _1411_ _0988_ _0989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2677_ _0937_ _0940_ _0941_ _0223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1628_ _1235_ _1245_ _1246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2325__A2 _0658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1559_ u1.timer\[27\] _1177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3229_ u1.row_col_select\[5\] clknet_leaf_21_clock net199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2089__A1 u0.cmd\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1836__A1 _0301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2261__A1 _0565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3045__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2541__I _0820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3195__CLK clknet_leaf_6_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2564__A2 _0852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2316__A2 _0630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1827__A1 _0299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2863__D control_trigger vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2252__A1 _1095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2451__I _1085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2600_ u1.row_sel\[1\] _0878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2531_ _0820_ _0833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2462_ _1085_ _0761_ _0754_ _0778_ _0779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__3282__I net98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2393_ _0708_ _0710_ _0718_ _0162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3014_ _0156_ clknet_leaf_37_clock u1.ordering_timer\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3068__CLK clknet_leaf_7_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2491__B2 _0565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2243__A1 _1062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2905__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2729_ _0281_ _1322_ _0974_ _0978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA_input52_I spi_data[20] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1705__I _1321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2085__I1 u1.ordering_complete\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2271__I _0610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2858__D u0.cmd\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1899__I1 _0345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3210__CLK clknet_leaf_36_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2928__CLK clknet_leaf_24_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1962_ _0392_ _0400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3277__I net108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1893_ u0.cmd\[19\] _0349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2514_ _0517_ _0818_ _0821_ spi_data_crossing\[1\].data_sync _0823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2445_ _1046_ _0763_ _0764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2000__I1 _0345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2376_ _1096_ _0703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3233__CLK clknet_leaf_22_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2455__A1 _0769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2058__I1 u1.ordering_complete\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2230_ _1102_ _1106_ _0572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2161_ _0529_ _0530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2092_ _1097_ _0455_ _0484_ _0095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_19_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2994_ _0136_ clknet_leaf_20_clock u1.row_col_select\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2461__A4 _0747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3106__CLK clknet_leaf_24_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1945_ u0.cmd\[14\] _0387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1876_ _0317_ _0333_ u1.col_sel\[2\] _0337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2221__I1 u1.row_col_select\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1724__A3 _1335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2428_ _0583_ u1.ordering_timer\[18\] _0723_ _0748_ _0749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_28_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2359_ _0670_ _0686_ _0688_ _0689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input15_I la_data_in[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1660__A2 _1277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3129__CLK clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1730_ _1164_ u1.ccr0\[25\] u1.ccr0\[24\] _1166_ _1346_ _1347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_11_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1784__B _1400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1661_ _1187_ _1222_ _1278_ _1279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1592_ _1207_ u1.ccr1\[0\] u1.ccr1\[1\] _1209_ _1210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3262_ clknet_leaf_12_clock net81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2213_ _0367_ u1.row_col_select\[5\] _0558_ _0560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3193_ _0263_ clknet_leaf_17_clock u1.ccr0\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1803__I _1327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input7_I la_data_in[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2144_ _0518_ _0113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2075_ _0474_ _1112_ _0470_ _0475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2977_ _0119_ clknet_leaf_17_clock u1.col_limit\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1928_ _0375_ _0040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1859_ u1.col_sel\[0\] _0321_ u1.col_sel\[1\] _0318_ _0322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_33_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1914__S _0354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2830__A1 net14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2649__A1 _1277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2900_ _0042_ clknet_leaf_25_clock u1.ccr0\[26\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1624__A2 _1236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2831_ _1039_ _0279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2762_ _1167_ _0998_ _0999_ _0934_ _0250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3285__I net101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1713_ _1327_ _1328_ _1329_ u1.timer\[22\] _1330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2693_ _1250_ _0951_ _0953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2188__I0 _0365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1644_ u1.timer\[12\] _1262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1575_ u1.timer\[7\] _1193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3245_ u0.mem_write_n\[1\] clknet_leaf_11_clock net183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3176_ net61 net72 spi_data_crossing\[29\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2127_ u0.cmd\[11\] _0507_ _0508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_2058_ _0462_ u1.ordering_complete\[3\] _0460_ _0463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2179__I0 _0513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output169_I net169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1551__A1 u1.ccr1\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2803__A1 _0468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2961__CLK clknet_leaf_33_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1790__A1 _1206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput81 net81 clock_out[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput92 net92 col_select_right[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__1542__B2 _1160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3030_ _0172_ clknet_leaf_30_clock u1.ordering_timer\[26\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2814_ _1296_ _1025_ _1030_ _0271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2745_ _0983_ _0987_ _0988_ _0244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_11_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2676_ u1.timer\[0\] u1.timer\[1\] u1.timer\[3\] u1.timer\[2\] _0941_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1627_ _1238_ _1244_ _1245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1558_ u1.ccr1\[27\] _1176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1489_ u1.ordering_timer\[11\] _1104_ u1.ordering_timer\[10\] _1113_ _1114_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3228_ u1.row_col_select\[4\] clknet_leaf_21_clock net198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2834__CLK clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2089__A2 _0478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1836__A2 _0305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3159_ spi_data_crossing\[20\].A clknet_leaf_8_clock spi_data_crossing\[20\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2984__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1901__I u0.cmd\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2530_ _0817_ _0832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2461_ _1064_ _0729_ _0777_ _0747_ _0778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__2857__CLK clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1515__A1 u1.ordering_timer\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2392_ _0329_ _0717_ _0718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3013_ _0155_ clknet_leaf_0_clock u1.ordering_timer\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2491__A2 _0709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1967__B _0403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2728_ _0281_ _0976_ _0977_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1754__A1 _1364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2659_ _1187_ _0926_ _0927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input45_I spi_data[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3125__D spi_data_crossing\[3\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3012__CLK clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3162__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1631__I u1.ccr1\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2473__A2 _0716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1961_ u0.cmd\[2\] _0399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1892_ _0347_ _0348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1984__A1 _1247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2513_ _0822_ _0178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2444_ _0754_ _0750_ _0763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2375_ _0702_ _0160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3035__CLK clknet_leaf_30_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3185__CLK clknet_leaf_36_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1917__S _0354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1451__I u1.ordering_timer\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2455__A2 _0755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1966__A1 _0402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3058__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2391__A1 _0711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2160_ _0528_ _0529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2694__A2 _0951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2091_ u0.cmd\[15\] _0478_ _0484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2993_ _0135_ clknet_leaf_22_clock u1.inverter_select\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1944_ _1357_ _0378_ _0386_ _0045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_37_clock_I clknet_2_0__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1875_ _0317_ u1.col_sel\[2\] _0333_ _0336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_30_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2427_ _0747_ _0748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2358_ u1.ordering_complete\[12\] _0687_ _0688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2289_ u1.ordering_timer\[0\] u1.ordering_timer\[1\] u1.ordering_timer\[3\] u1.ordering_timer\[2\]
+ _0627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_38_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3200__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1446__I u1.ordering_timer\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2373__A1 _0670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2918__CLK clknet_leaf_34_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2226__B _1137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1660_ _1246_ _1277_ _1278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1591_ _1208_ _1209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3261_ clknet_leaf_12_clock net80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2116__A1 u0.cmd\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2212_ _0559_ _0140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3192_ _0262_ clknet_leaf_16_clock u1.ccr0\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2143_ _0517_ u1.row_limit\[1\] _0515_ _0518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2187__I _0539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2074_ u0.cmd\[8\] _0474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3223__CLK clknet_leaf_22_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2976_ _0118_ clknet_leaf_14_clock u1.row_limit\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1927_ u1.ccr0\[24\] _0374_ _0358_ _0375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1858_ u1.col_limit\[0\] _0321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1789_ _1289_ _1280_ _1283_ _1287_ _1406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__2658__A2 _0918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2097__I _0488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1930__S _0358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1904__I _0352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1857__B1 u1.col_sel\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2890__CLK clknet_leaf_23_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2649__A2 _0916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3246__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2735__I _0933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2821__A2 _1015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2830_ net14 net32 _1039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_32_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2761_ u1.timer\[30\] _0996_ _1413_ _0993_ _0999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1712_ u1.ccr0\[22\] _1329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2692_ _0946_ _0951_ _0952_ _0227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1643_ u1.ccr1\[12\] _1261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_0_clock_I clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1574_ u1.ccr1\[6\] _1189_ u1.ccr1\[5\] _1191_ _1192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3244_ u0.mem_write_n\[0\] clknet_leaf_11_clock net182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3175_ spi_data_crossing\[28\].A clknet_leaf_11_clock spi_data_crossing\[28\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2126_ _0486_ _0507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_2057_ _0402_ _0462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2959_ _0101_ clknet_leaf_33_clock u1.ordering_complete\[21\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3119__CLK clknet_leaf_38_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_6_clock_I clknet_2_1__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1551__A2 _1167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2500__A1 u1.ordering_timer\[27\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2803__A2 _1021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1917__I1 _0367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput82 net82 clock_out[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput93 net93 col_select_right[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_23_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3296__I net162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2813_ u0.cmd\[10\] _1029_ _1030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2558__A1 u0.cmd\[18\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2744_ u1.timer\[24\] _1327_ _0286_ _0981_ _0988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_9_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2675_ _1214_ _0938_ _0940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1626_ _1241_ _1242_ _1243_ _1244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_28_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1557_ _1172_ _1174_ _1175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1533__A2 u0.cmd\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2730__A1 _0968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1488_ u1.ordering_complete\[10\] _1113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3227_ u1.row_col_select\[3\] clknet_leaf_21_clock net197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3158_ net52 net72 spi_data_crossing\[20\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2109_ _0464_ u1.ordering_complete\[20\] _0496_ _0497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3089_ _0223_ clknet_leaf_5_clock u1.timer\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2721__A1 _1279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2721__B2 _0283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1454__I u1.ordering_complete\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3091__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2234__B _1108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1763__A2 _1290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2460_ _0703_ _0698_ _0776_ _0722_ _0777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_29_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2391_ _0711_ _0713_ _0715_ _0716_ _0717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2712__A1 _1254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3012_ _0154_ clknet_leaf_0_clock u1.ordering_timer\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2727_ _0968_ _0975_ _0976_ _0238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2658_ _1246_ _0918_ _0925_ _0926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2589_ _0868_ _0208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1609_ _1225_ u1.timer\[23\] _1226_ u1.timer\[22\] _1227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1506__A2 u1.ordering_complete\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2703__A1 _0958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input38_I la_oenb[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2951__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1993__A2 _0416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1960_ _0397_ _0398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1891_ u0.cmd\[17\] _0347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2512_ _0513_ _0818_ _0821_ spi_data_crossing\[0\].data_sync _0822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3226__D u1.row_col_select\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2974__CLK clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2443_ _0602_ _0762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2374_ _0698_ _0682_ _0691_ _0701_ _0702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_33_clock_I clknet_2_2__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2449__B1 _0762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2847__CLK clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1966__A2 _0400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2215__I0 _0369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2997__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1907__I _0353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2090_ _1098_ _0455_ _0483_ _0094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_46_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2446__A3 _0750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2992_ _0134_ clknet_leaf_22_clock u1.inverter_select\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1943_ _0385_ _0383_ _0386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1874_ _0331_ _0335_ _0026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2206__I0 _0360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3002__CLK clknet_leaf_22_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2426_ u1.ordering_timer\[21\] u1.ordering_timer\[20\] _0747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3152__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2134__A2 _0490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2357_ _0629_ _0687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2288_ _0625_ _0626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2383__I _0624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1462__I u1.ordering_timer\[26\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1884__A1 _0311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2428__A3 _0723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3025__CLK clknet_leaf_32_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3175__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1590_ u1.timer\[1\] _1208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3260_ clknet_leaf_12_clock net79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2116__A2 _0493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2211_ _0365_ u1.row_col_select\[4\] _0558_ _0559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3191_ _0261_ clknet_leaf_16_clock u1.ccr0\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2142_ _0457_ _0517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2073_ _0473_ _0087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3299__I net165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2975_ _0117_ clknet_leaf_15_clock u1.row_limit\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1926_ u0.cmd\[8\] _0374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1857_ _0317_ _0318_ u1.col_sel\[2\] _0319_ _0320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1547__I u1.timer\[24\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1788_ _1256_ _1257_ _1258_ _1404_ _1405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2355__A2 _0675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2107__A2 _0489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2409_ _0329_ _0732_ _0733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input20_I la_data_in[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output107_I net107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3048__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_2_clock_I clknet_2_0__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3198__CLK clknet_leaf_6_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2346__A2 _0665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1554__B1 u1.ccr1\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2288__I _0625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1920__I _0353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1609__B2 u1.timer\[22\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2282__A1 _0611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2760_ _0996_ _0995_ _0998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1711_ u1.ccr0\[23\] _1328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2691_ _1289_ _0948_ _0952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1642_ _1255_ _1259_ _1260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1573_ _1190_ _1191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3312_ net209 net215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3243_ u0.cmd\[25\] clknet_leaf_11_clock net171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3234__D u0.cmd\[16\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3174_ net60 net72 spi_data_crossing\[28\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2125_ u1.ordering_complete\[27\] _0506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_2056_ _0461_ _0082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2273__A1 _1138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_2_2__f_clock_I clknet_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2908__CLK clknet_leaf_15_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2958_ _0100_ clknet_leaf_34_clock u1.ordering_complete\[20\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1909_ _1320_ _0359_ _0362_ _0034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2889_ u1.u1.impulse_gen\[0\] clknet_leaf_17_clock u1.u1.impulse_gen\[1\] vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input68_I spi_data[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2264__A1 _1138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1790__A3 _1214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput83 net83 col_select_left[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput94 net94 col_select_right[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__3213__CLK clknet_leaf_36_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2812_ _1011_ _1029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2743_ _0285_ _0985_ u1.timer\[24\] _0987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2674_ _0937_ _0938_ _0939_ _0222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1625_ u1.ccr1\[16\] _1237_ _1243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2430__B _0750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1556_ u1.ccr1\[29\] _1168_ u1.ccr1\[28\] _1173_ _1174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1533__A3 _1042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1487_ u1.ordering_complete\[8\] _1112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3226_ u1.row_col_select\[2\] clknet_leaf_21_clock net196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_2_3__f_clock clknet_0_clock clknet_2_3__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3157_ spi_data_crossing\[19\].A clknet_leaf_8_clock spi_data_crossing\[19\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2494__A1 u1.ordering_timer\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2108_ _0487_ _0496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_42_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3088_ _0222_ clknet_leaf_5_clock u1.timer\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2039_ u0.cmd\[16\] _0447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2880__CLK clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_28_clock_I clknet_2_2__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3139__D spi_data_crossing\[10\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output174_I net174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3236__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1735__I u1.ccr0\[31\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2021__I1 _0374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2485__A1 u1.ordering_complete\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2237__A1 _1187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1645__I u1.ccr1\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2390_ _0624_ _0716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2476__A1 u1.ordering_timer\[27\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3011_ _0153_ clknet_leaf_0_clock u1.ordering_timer\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2228__B2 _1129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2228__A1 _1132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3109__CLK clknet_leaf_24_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2726_ _1321_ _0282_ u1.timer\[16\] _0970_ _0976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2657_ _0919_ _1234_ _1235_ _0923_ _0924_ _0925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__1555__I u1.timer\[28\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1608_ u1.ccr1\[22\] _1226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2588_ u0.cmd\[30\] _0864_ _0865_ spi_data_crossing\[30\].data_sync _0868_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1539_ _1158_ _0011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3209_ _0001_ clknet_leaf_38_clock net161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output99_I net99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2458__A1 _0648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1681__A2 _1296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2630__A1 _0891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1890_ u0.cmd\[16\] _0346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2511_ _0820_ _0821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2442_ u1.ordering_timer\[23\] _0761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2373_ _0670_ _0699_ _0700_ _0701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2697__A1 _0951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3081__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2621__A1 _0890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2709_ _0958_ _0963_ _0964_ _0232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_input50_I spi_data[19] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2688__A1 _0946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output137_I net137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2612__A1 _0875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1923__I u0.cmd\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2991_ _0133_ clknet_leaf_21_clock u1.inverter_select\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1942_ u0.cmd\[13\] _0385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1873_ _0317_ _0333_ _0335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2941__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2206__I1 u1.row_col_select\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3237__D u0.cmd\[19\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2425_ u1.ordering_timer\[20\] _0737_ _0746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2356_ _0684_ _0685_ _0686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2287_ _0624_ _0625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2964__CLK clknet_leaf_33_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2015__S _0427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2364__A3 _0665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2210_ _0552_ _0558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3190_ _0260_ clknet_leaf_38_clock net151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1875__A2 u1.col_sel\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2141_ _0516_ _0112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2072_ _0472_ u1.ordering_complete\[7\] _0470_ _0473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2824__A1 u0.cmd\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2974_ _0116_ clknet_leaf_14_clock u1.row_limit\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2588__B1 _0865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1925_ _1328_ _0359_ _0373_ _0039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2052__A2 _0453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1856_ u1.col_limit\[2\] _0319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1787_ _1311_ _1404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2355__A3 _0677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2837__CLK clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2408_ _0711_ _0730_ _0731_ _0716_ _0732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_44_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2339_ u1.ordering_timer\[10\] _0665_ _0671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input13_I la_data_in[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2394__I _0625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2987__CLK clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1554__B2 _1167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1554__A1 u1.ccr1\[31\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1857__A2 _0318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2806__A1 _0372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1490__B1 _1111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3142__CLK net72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1710_ u1.timer\[23\] _1327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2690_ _0950_ _0951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1641_ u1.ccr1\[15\] _1256_ u1.ccr1\[14\] _1257_ u1.ccr1\[13\] _1258_ _1259_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3311_ net208 net214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1572_ u1.timer\[5\] _1190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3242_ u0.cmd\[24\] clknet_leaf_11_clock net170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3173_ spi_data_crossing\[27\].A clknet_leaf_10_clock spi_data_crossing\[27\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input5_I la_data_in[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2124_ _0504_ _0500_ _0505_ _0106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2055_ _0459_ u1.ordering_complete\[2\] _0460_ _0461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2957_ _0099_ clknet_leaf_33_clock u1.ordering_complete\[19\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2888_ u1.ccr1_flag clknet_leaf_17_clock u1.u1.impulse_gen\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1908_ _0360_ _0361_ _0362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1839_ _0304_ _1153_ _0298_ _0020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1784__A1 _1292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_24_clock_I clknet_2_3__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3015__CLK clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2500__A3 _0769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3165__CLK clknet_leaf_10_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1775__A1 _1337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput84 net84 col_select_left[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput73 net73 clock_out[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput95 net95 data_out_left[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_27_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2811_ _1028_ _0270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2742_ _0285_ _0985_ _0986_ _0982_ _0243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_9_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2673_ _1206_ _1208_ _1203_ _0939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1624_ u1.ccr1\[17\] _1236_ _1242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1518__A1 _1132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3038__CLK clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1555_ u1.timer\[28\] _1173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2730__A3 _0978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3225_ u1.row_col_select\[1\] clknet_leaf_21_clock net195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1486_ u1.ordering_timer\[8\] _1111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_45_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3156_ net50 net72 spi_data_crossing\[19\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3188__CLK clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2494__A2 _0791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3087_ _0221_ clknet_leaf_5_clock u1.timer\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2107_ _1058_ _0489_ _0495_ _0099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2038_ _0446_ _0079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2113__S _0496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output167_I net167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2485__A2 _0720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2237__A2 _1235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1996__A1 _0389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1748__A1 _1363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1748__B2 _1364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2796__I0 u1.ccr0\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1926__I u0.cmd\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2757__I u1.timer\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3010_ _0152_ clknet_leaf_0_clock u1.ordering_timer\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2228__A2 _0568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1739__A1 _1348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2725_ _1322_ _0974_ _0975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2656_ u1.ccr1\[23\] _1228_ _1227_ _0924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1607_ u1.ccr1\[23\] _1225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2587_ _0867_ _0207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2164__A1 _0321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1538_ u0.run_state\[3\] u0.run_state\[4\] _1158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1911__A1 _0363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1469_ _1093_ u1.ordering_complete\[27\] _1087_ u1.ordering_complete\[26\] _1094_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__2667__I _0934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3208_ _0278_ clknet_leaf_38_clock net158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3139_ spi_data_crossing\[10\].A clknet_leaf_2_clock spi_data_crossing\[10\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1978__A1 _0372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3203__CLK clknet_leaf_7_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1969__A1 _0404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2510_ _0819_ _0820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2441_ _0760_ _0168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2372_ u1.ordering_complete\[14\] _0687_ _0700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2870__CLK clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2449__A2 _0755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3226__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2708_ _1311_ _0961_ _0964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2639_ _0906_ _1270_ _0907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input43_I spi_data[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2679__A2 _0941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2893__CLK clknet_leaf_26_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3249__CLK clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2990_ _0132_ clknet_leaf_22_clock u1.inverter_select\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1941_ _1358_ _0378_ _0384_ _0044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1872_ _0331_ _0333_ _0334_ _0025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2211__S _0558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2424_ _0745_ _0166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2355_ u1.ordering_timer\[12\] _0675_ _0677_ _0685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_9_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2010__I _0422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2286_ _0600_ _0624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2358__A1 u1.ordering_complete\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2597__A1 _0309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_19_clock_I clknet_2_3__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2349__A1 _0670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2364__A4 _0692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2031__S _0438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3071__CLK clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2140_ _0513_ u1.row_limit\[0\] _0515_ _0516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2765__I net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2071_ u0.cmd\[7\] _0472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2973_ _0115_ clknet_leaf_14_clock u1.row_limit\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2588__A1 u0.cmd\[30\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2588__B2 spi_data_crossing\[30\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1924_ _0372_ _0370_ _0373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1855_ u1.col_limit\[1\] _0318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2005__I _0426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1786_ _1402_ _1144_ _1403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1563__A2 _1180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2512__A1 _0513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2407_ u1.ordering_complete\[18\] _0725_ _0731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2512__B2 spi_data_crossing\[0\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2338_ _0610_ _0670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2269_ _0609_ _0147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_20_clock_I clknet_2_3__leaf_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1955__S _0394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3094__CLK clknet_leaf_4_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1554__A2 _1171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2503__A1 _0603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2931__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2806__A2 _1021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1490__A1 _1109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1490__B2 _1112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1929__I u0.cmd\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3068__D _0023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1640_ u1.timer\[13\] _1258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1571_ _1188_ _1189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3310_ net207 net213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3241_ u0.cmd\[23\] clknet_leaf_10_clock net169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3172_ net59 net72 spi_data_crossing\[27\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2123_ u0.cmd\[10\] _0493_ _0505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2054_ _0452_ _0460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_19_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1481__B2 u1.ordering_complete\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2956_ _0098_ clknet_leaf_34_clock u1.ordering_complete\[18\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2887_ _0021_ clknet_leaf_12_clock u0.mem_write_n\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1907_ _0353_ _0361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1838_ _0299_ _1160_ _0302_ _0305_ _0019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2033__I0 u1.ccr1\[29\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1769_ _1375_ _1381_ _1383_ _1384_ _1385_ _1386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_1_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2954__CLK clknet_leaf_34_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1839__A3 _0298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2500__A4 _0784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2024__I0 u1.ccr1\[25\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1527__A2 _1044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2724__A1 _0968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput85 net85 col_select_left[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput74 net74 clock_out[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput96 net96 data_out_left[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_49_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2810_ u1.ccr0\[9\] _0376_ _1013_ _1028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2741_ _0285_ _0985_ _0986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2672_ _1364_ _1363_ _1204_ _0938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2977__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1623_ _1239_ _1240_ _1241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1554_ u1.ccr1\[31\] _1171_ u1.ccr1\[30\] _1167_ _1172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_28_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1485_ u1.ordering_complete\[9\] _1110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3224_ u1.row_col_select\[0\] clknet_leaf_21_clock net194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

